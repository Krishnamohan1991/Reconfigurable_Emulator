module FPGA_testbench();
//reg clk,reset,prgm_b,cb_prgm_b;

integer input_file;

reg [767:0] CB_config_stream ;
reg [1183:0] CLB_config_stream;
reg [191:0] IO_config_stream;
reg [6912:0] SB_config_stream;


reg [767:0] CB_config_stream_final ;
reg [1183:0] CLB_config_stream_final;
reg [191:0] IO_config_stream_final;
reg [6912:0] SB_config_stream_final;
//reg [3071:0] SB_config_stream;


//reg [1535:0] SB_config_stream;
//reg [1535:0] SB_config_stream_2;

//reg [3071:0] SB_config_stream_3;
wire cb_prgm_b_out,cb_prgm_b_out_1;
wire G0,G1,G2,G3,G4,G5,G6,G7;
integer i,k,l,m;


inout V00_0,V00_1,V00_2,V00_3,V00_4,V00_5,V00_6,V00_7,V01_0,V01_1,V01_2,V01_3,V01_4,V01_5,V01_6,V01_7,
	    V02_0,V02_1,V02_2,V02_3,V02_4,V02_5,V02_6,V02_7,V10_0,V10_1,V10_2,V10_3,V10_4,V10_5,V10_6,V10_7,
	    V11_0,V11_1,V11_2,V11_3,V11_4,V11_5,V11_6,V11_7,V12_0,V12_1,V12_2,V12_3,V12_4,V12_5,V12_6,V12_7,
            H00_0,H00_1,H00_2,H00_3,H00_4,H00_5,H00_6,H00_7,H01_0,H01_1,H01_2,H01_3,H01_4,H01_5,H01_6,H01_7,
	    H10_0,H10_1,H10_2,H10_3,H10_4,H10_5,H10_6,H10_7,H11_0,H11_1,H11_2,H11_3,H11_4,H11_5,H11_6,H11_7,
	    H20_0,H20_1,H20_2,H20_3,H20_4,H20_5,H20_6,H20_7,H21_0,H21_1,H21_2,H21_3,H21_4,H21_5,H21_6,H21_7;



 reg H000,H001,H002,H003,H004,H005,H006,H007,H010,H011,H012,H013,H014,H015,H016,H017,
	   H100,H101,H102,H103,H104,H105,H106,H107,H110,H111,H112,H113,H114,H115,H116,H117,
	   H200,H201,H202,H203,H204,H205,H206,H207,H210,H211,H212,H213,H214,H215,H216,H217;
 
 reg V000,V001,V002,V003,V004,V005,V006,V007,V010,V011,V012,V013,V014,V015,V016,V017,
	    V020,V021,V022,V023,V024,V025,V026,V027,V100,V101,V102,V103,V104,V105,V106,V107,
	    V110,V111,V112,V113,V114,V115,V116,V117,V120,V121,V122,V123,V124,V125,V126,V127;
 
value v0(.in(V000),.out(V00_0));         value v24(.in(V100),.out(V10_0));
value v1(.in(V001),.out(V00_1));         value v25(.in(V101),.out(V10_1));
value v2(.in(V002),.out(V00_2));         value v26(.in(V102),.out(V10_2));
value v3(.in(V003),.out(V00_3));         value v27(.in(V103),.out(V10_3));
value v4(.in(V004),.out(V00_4));         value v28(.in(V104),.out(V10_4));
value v5(.in(V005),.out(V00_5));         value v29(.in(V105),.out(V10_5));
value v6(.in(V006),.out(V00_6));         value v30(.in(V106),.out(V10_6));
value v7(.in(V007),.out(V00_7));         value v31(.in(V107),.out(V10_7));
value v8(.in(V010),.out(V01_0));         //value v32(.in(V110),.out(V11_0)); 
value v9(.in(V011),.out(V01_1));         value v33(.in(V111),.out(V11_1)); 
value v10(.in(V012),.out(V01_2));        value v34(.in(V112),.out(V11_2));
value v11(.in(V013),.out(V01_3));        value v35(.in(V113),.out(V11_3)); 
value v12(.in(V014),.out(V01_4));        value v36(.in(V114),.out(V11_4)); 
value v13(.in(V015),.out(V01_5));        value v37(.in(V115),.out(V11_5)); 
value v14(.in(V016),.out(V01_6));        value v38(.in(V116),.out(V11_6)); 
value v15(.in(V017),.out(V01_7));        value v39(.in(V117),.out(V11_7));
value v16(.in(V020),.out(V02_0));        value v40(.in(V120),.out(V12_0));
value v17(.in(V021),.out(V02_1));        value v41(.in(V121),.out(V12_1));
value v18(.in(V022),.out(V02_2));        value v42(.in(V122),.out(V12_2));
value v19(.in(V023),.out(V02_3));        value v43(.in(V123),.out(V12_3));
value v20(.in(V024),.out(V02_4));        value v44(.in(V124),.out(V12_4));
value v21(.in(V025),.out(V02_5));        value v45(.in(V125),.out(V12_5));
value v22(.in(V026),.out(V02_6));        value v46(.in(V126),.out(V12_6));
value v23(.in(V027),.out(V02_7));        value v47(.in(V127),.out(V12_7));

value H0(.in(H000),.out(H00_0));         value H24(.in(H100),.out(H10_0));
value H1(.in(H001),.out(H00_1));         value H25(.in(H101),.out(H10_1));
value H2(.in(H002),.out(H00_2));         value H26(.in(H102),.out(H10_2));
value H3(.in(H003),.out(H00_3));         value H27(.in(H103),.out(H10_3));
value H4(.in(H004),.out(H00_4));         value H28(.in(H104),.out(H10_4));
value H5(.in(H005),.out(H00_5));         value H29(.in(H105),.out(H10_5));
value H6(.in(H006),.out(H00_6));         value H30(.in(H106),.out(H10_6));
value H7(.in(H007),.out(H00_7));         value H31(.in(H107),.out(H10_7));
value H8(.in(H010),.out(H01_0));         value H32(.in(H110),.out(H11_0));
value H9(.in(H011),.out(H01_1));         value H33(.in(H111),.out(H11_1));
value H10(.in(H012),.out(H01_2));        value H34(.in(H112),.out(H11_2));
value H11(.in(H013),.out(H01_3));        value H35(.in(H113),.out(H11_3));
value H12(.in(H014),.out(H01_4));        value H36(.in(H114),.out(H11_4));
value H13(.in(H015),.out(H01_5));        value H37(.in(H115),.out(H11_5));
value H14(.in(H016),.out(H01_6));        value H38(.in(H116),.out(H11_6));
value H15(.in(H017),.out(H01_7));        value H39(.in(H117),.out(H11_7));
value H16(.in(H020),.out(H02_0));        value H40(.in(H120),.out(H12_0));
value H17(.in(H021),.out(H02_1));        value H41(.in(H121),.out(H12_1));
value H18(.in(H022),.out(H02_2));        value H42(.in(H122),.out(H12_2));
value H19(.in(H023),.out(H02_3));        value H43(.in(H123),.out(H12_3));
value H20(.in(H024),.out(H02_4));        value H44(.in(H124),.out(H12_4));
value H21(.in(H025),.out(H02_5));        value H45(.in(H125),.out(H12_5));
value H22(.in(H026),.out(H02_6));        value H46(.in(H126),.out(H12_6));
value H23(.in(H027),.out(H02_7));        value H47(.in(H127),.out(H12_7));


     

reg clk,reset,prgm_b,CLB_prgm_b,cb_prgm_b,sb_prgm_b,bit_in_CLB,bit_in_CB,bit_in_SB,bit_in_SB_2,sb_prgm_b_in,
cb_prgm_b_in,CLB_prgm_b_in,sb_prgm_b_2,io_prgm_b_in,bit_in_IO,io_prgm_b;

integer CB_count,SB_count,SB_count_2,CLB_count,CLB_counter,CB_counter,SB_counter,SB_counter_2,IO_counter,IO_count;


FPGA FPGA1(.V00_0(V00_0),.V00_1(V00_1),.V00_2(V00_2),.V00_3(V00_3),
.V00_4(V00_4),.V00_5(V00_5),.V00_6(V00_6),.V00_7(V00_7),.V01_0(V01_0),
.V01_1(V01_1),.V01_2(V01_2),.V01_3(V01_3),.V01_4(V01_4),.V01_5(V01_5),
.V01_6(V01_6),.V01_7(V01_7),.V02_0(V02_0),.V02_1(V02_1),.V02_2(V02_2),
.V02_3(V02_3),.V02_4(V02_4),.V02_5(V02_5),.V02_6(V02_6),.V02_7(V02_7),
.V10_0(V10_0),.V10_1(V10_1),.V10_2(V10_2),.V10_3(V10_3),.V10_4(V10_4),
.V10_5(V10_5),.V10_6(V10_6),.V10_7(V10_7),.V11_0(V11_0),.V11_1(V11_1),
.V11_2(V11_2),.V11_3(V11_3),.V11_4(V11_4),.V11_5(V11_5),.V11_6(V11_6),
.V11_7(V11_7),.V12_0(V12_0),.V12_1(V12_1),.V12_2(V12_2),.V12_3(V12_3),
.V12_4(V12_4),.V12_5(V12_5),.V12_6(V12_6),.V12_7(V12_7),.H00_0(H00_0),
.H00_1(H00_1),.H00_2(H00_2),.H00_3(H00_3),.H00_4(H00_4),.H00_5(H00_5),
.H00_6(H00_6),.H00_7(H00_7),.H01_0(H01_0),.H01_1(H01_1),.H01_2(H01_2),
.H01_3(H01_3),.H01_4(H01_4),.H01_5(H01_5),.H01_6(H01_6),.H01_7(H01_7),
.H10_0(H10_0),.H10_1(H10_1),.H10_2(H10_2),.H10_3(H10_3),.H10_4(H10_4),
.H10_5(H10_5),.H10_6(H10_6),.H10_7(H10_7),.H11_0(H11_0),.H11_1(H11_1),
.H11_2(H11_2),.H11_3(H11_3),.H11_4(H11_4),.H11_5(H11_5),.H11_6(H11_6),
.H11_7(H11_7),.H20_0(H20_0),.H20_1(H20_1),.H20_2(H20_2),.H20_3(H20_3),
.H20_4(H20_4),.H20_5(H20_5),.H20_6(H20_6),.H20_7(H20_7),.H21_0(H21_0),
.H21_1(H21_1),.H21_2(H21_2),.clk(clk),.reset(reset),.prgm_b(prgm_b),
.CLB_prgm_b(CLB_prgm_b),.cb_prgm_b(cb_prgm_b),.sb_prgm_b(sb_prgm_b),
.sb_prgm_b_2(sb_prgm_b_2),.bit_in_CLB(bit_in_CLB),.bit_in_CB(bit_in_CB),
.sb_prgm_b_in(sb_prgm_b_in),.cb_prgm_b_in(cb_prgm_b_in),.CLB_prgm_b_in(CLB_prgm_b_in),
.bit_in_SB(bit_in_SB),.bit_in_SB_2(bit_in_SB_2),.io_prgm_b(io_prgm_b),.bit_in_IO(bit_in_IO),.io_prgm_b_in(io_prgm_b_in)); 

//For all bit-streams the bits are arranged in the decreasing order of their coordinate positions. eg. The bits belonging to the first CLB CLB_00 will be placed at the end of the CLB bitstream

initial begin
//input_file=$fopen("/home/krishna/Downloads/DEV_Git/conf_bit_stream.txt","r");
clk = 1'b0;
 reset=1'b0;
 
 prgm_b=1'b1;   //indicates start of bit_stream----active low
 cb_prgm_b=1'b0;
 cb_prgm_b_in=1'b0;
 sb_prgm_b=1'b0;
 sb_prgm_b_in=1'b0;
 sb_prgm_b_2=1'b0;
 CLB_prgm_b=1'b0;
 io_prgm_b_in=1'b0;
 io_prgm_b=1'b0;

 fork
/*
 #1 while(!$feof(input_file))
	begin
	CB_config_stream_final=$fscanf(input_file,"%b\n",CB_config_stream);
	SB_config_stream_final=$fscanf(input_file,"%b\n",SB_config_stream);
	CLB_config_stream_final=$fscanf(input_file,"%b\n",CLB_config_stream);
	IO_config_stream_final=$fscanf(input_file,"%b\n",IO_config_stream);
	end
	$fclose(input_file);
*/
 #1 reset=1'b1;
 #1 prgm_b=1'b0;
 #1 cb_prgm_b=1'b1;
 #1 cb_prgm_b_in=1'b1;
 #1 sb_prgm_b=1'b1;
 #1 sb_prgm_b_2=1'b1;
 #1 sb_prgm_b_in=1'b1;
 #1 CLB_prgm_b=1'b1;
 #1 CLB_prgm_b_in=1'b1;
 #1 io_prgm_b_in=1'b1;
 #1 io_prgm_b=1'b1;

 #1 CB_counter=0;CB_count=0;
 #1 CLB_counter=0;CLB_count=0;
 #1 SB_counter=0;SB_count=0;
 #1 SB_counter_2=0;SB_count_2=0;
 #1 IO_counter=0;IO_count=0;
 #1 reset=1'b1;
 #2 reset=1'b0;

 join
end

initial begin
//for(i=0;i<=6074;i++)
//begin

forever #5 clk=!clk;

end

initial
begin

CB_config_stream[767:0]= 768'b000000000000000000000000000000000000000000000000100000010000001000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000010000001000000100000010000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
SB_config_stream[6911:0]= 6912'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000010000000000000000010000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
CLB_config_stream[1183:0]= 1184'b00000000000000000000100000000000000000000000000000000000010000000000000000010000100101010010111100000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000001000000000000000000000000010001000011110000000000000000000000001000100001111000000000000000;
IO_config_stream[191:0]=192'b000000000000000010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110100000000000000000000000000000000000001111111110100000;

for(i=0;i<6912;i=i+1)
SB_config_stream_final[i]=SB_config_stream[i];

for(k=0;k<1184;k=k+1)
CLB_config_stream_final[k]=CLB_config_stream[k];

for(l=0;l<768;l=l+1)
CB_config_stream_final[l]=CB_config_stream[l];

for(m=0;m<192;m=m+1)
IO_config_stream_final[m]=IO_config_stream[m];


end

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && cb_prgm_b!=1'b0) begin

	
	
    if((CB_counter == 49) && cb_prgm_b!=1'b0) //(no of bits required for one CB) + 1= 48+1=49
	begin
	    
		CB_count=CB_count+1;
		
		CB_counter=0;
		if(CB_count==16)
		begin
			
			cb_prgm_b=1'b0;
           // prgm_b=1'b1;
			
		end
	end 
	bit_in_CB <= CB_config_stream_final[0];
	CB_config_stream_final <=CB_config_stream_final>>1;
	CB_counter=CB_counter+1;//if endsj
end 

end //always block ends


always@(posedge clk or posedge reset)
begin 

	if(prgm_b!=1'b1 && sb_prgm_b!=1'b0) begin
	
		if((SB_counter == 769) && sb_prgm_b!=1'b0) //(no of bits required for one SB +1 = 769)
			begin
	    
			SB_count=SB_count+1;
			SB_counter=0;
			if(SB_count==9)
			begin
			
				sb_prgm_b=1'b0;
			//sb_prgm_b_in=1'b1;
			 prgm_b=1'b1;
			
			end
		end 
	bit_in_SB <= SB_config_stream_final[0];
	SB_config_stream_final <=SB_config_stream_final>>1;
	SB_counter=SB_counter+1;//if endsj
	end 

end //always block ends
/*
always@(posedge clk or posedge reset)
begin 

	if(prgm_b!=1'b1 && sb_prgm_b_2!=1'b0) begin
	
		if((SB_counter_2 == 769) && sb_prgm_b_2!=1'b0) //(no of bits required for one SB +1 = 769)
			begin
	    
			SB_count_2=SB_count_2+1;
			SB_counter_2=0;
			if(SB_count_2==2)
			begin
			
				sb_prgm_b_2=1'b0;
			sb_prgm_b_in=1'b1;
			if(sb_prgm_b_2==1'b0)
			 	 prgm_b=1'b1;
			
			end
		end 
	bit_in_SB_2 <= SB_config_stream_2[0];
	SB_config_stream_2 <=SB_config_stream_2>>1;
	SB_counter_2=SB_counter_2+1;//if endsj
	end 

end //always block ends  

 */

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && CLB_prgm_b!=1'b0) 
begin

    if((CLB_counter == 297) && CLB_prgm_b!=1'b0) //(no of bits required for one CLB) + 1= 37+1=38  or (37 + (number of LUT -1))
	begin
	    
		CLB_count=CLB_count+1;
		
		CLB_counter=0;
		if(CLB_count==4)
		begin
			
			CLB_prgm_b=1'b0;
          
			
		end
	end 
	bit_in_CLB <= CLB_config_stream_final[0];
	CLB_config_stream_final <=CLB_config_stream_final>>1;
	CLB_counter=CLB_counter+1;//if endsj
end 

end //always block ends

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && io_prgm_b!=1'b0) 
begin	
	
    if((IO_counter == 17) && io_prgm_b!=1'b0) //(no of bits required for one IO block configuration + 1= 16+1=17
	begin
	    
		IO_count=IO_count+1;
		
		IO_counter=0;
		if(IO_count==12)
		begin
			
			io_prgm_b=1'b0;
           // prgm_b=1'b1;
			
		end
	end 
	bit_in_IO <= IO_config_stream_final[0];
	IO_config_stream_final <=IO_config_stream_final>>1;
	IO_counter=IO_counter+1;//if endsj
end 

end //always block ends

//end  

initial
	begin 
#600;               //time=5 seconds
V000=1;V001=1;V002=1;V003=1;//H05=1;H06=1;H07=1;H08=1;
H000=0;H001=1;H002=0;H003=1;
//V10=1;V11=1;
#800;
	//reset=1'b0;
V000=1;V001=1;V002=1;V003=1;//H05=1;H06=1;H07=1;H08=1;
H000=0;H001=1;H002=0;H003=1;
#800;
	//reset=1'b0;
V000=1;V001=1;V002=1;V003=1;//H05=1;H06=1;H07=1;H08=1;
H000=0;H001=1;H002=0;H003=1;
//V10=1;V11=1;
#86400 $finish;
end
initial begin
    $dumpfile("test.vcd");

    $dumpvars(0,FPGA_testbench);
    $timeformat(-9, 1, " ns", 6);
	$monitor("At prgm_b=%b reset=%b SB_count=%d",prgm_b,reset,SB_count);
end

//Stimulus

endmodule
