module FPGA_testbench();
//reg clk,reset,prgm_b,cb_prgm_b;

reg [767:0] CB_config_stream ;
reg [1183:0] CLB_config_stream;
reg [191:0] IO_config_stream;
reg [6912:0] SB_config_stream;


reg [767:0] CB_config_stream_final ;
reg [1183:0] CLB_config_stream_final;
reg [191:0] IO_config_stream_final;
reg [6912:0] SB_config_stream_final;
reg [3071:0]SB_config_stream_3;
reg [1535:0]SB_config_stream_2;
//reg [3071:0] SB_config_stream;


//reg [1535:0] SB_config_stream;
//reg [1535:0] SB_config_stream_2;

//reg [3071:0] SB_config_stream_3;
wire cb_prgm_b_out,cb_prgm_b_out_1;
wire G0,G1,G2,G3,G4,G5,G6,G7;
integer i;

inout V0_0,V0_1,V0_2,V0_3,V0_4,V0_5,V0_6,V0_7,V1_0,V1_1,V1_2,V1_3,V1_4,V1_5,V1_6,V1_7,
            H0_0,H0_1,H0_2,H0_3,H0_4,H0_5,H0_6,H0_7,H1_0,H1_1,H1_2,H1_3,H1_4,H1_5,H1_6,H1_7;
 reg H00,H01,H02,H03,H04,H05,H06,H07,V10,V11;
 reg V00,V01,V02,V03,V04;
/*
 value v1(.in(V00),.out(V0_0));  
 value v2(.in(V01),.out(V0_1));  
 value v3(.in(V02),.out(V0_2));  
 value v4(.in(V03),.out(V0_3)); 

value v5(.in(H00),.out(H0_0));  
 value v6(.in(H01),.out(H0_1));  
 value v7(.in(H02),.out(H0_2));  
 value v8(.in(H03),.out(H0_3)); */

 //value v5(.in(V10),.out(V1_0));  
 //value v6(.in(V11),.out(V1_1));  
 //value v7(.in(H07),.out(H0_6));  
 //value v8(.in(H08),.out(H0_7));          

reg clk,reset,prgm_b,CLB_prgm_b,cb_prgm_b,sb_prgm_b,bit_in_CLB,bit_in_CB,bit_in_SB,bit_in_SB_2,sb_prgm_b_in,cb_prgm_b_in,CLB_prgm_b_in,sb_prgm_b_2;

integer CB_count,SB_count,SB_count_2,CLB_count,CLB_counter,CB_counter,SB_counter,SB_counter_2;

FPGA FPGA1(.V0_0(V0_0),.V0_1(V0_1),.V0_2(V0_2),.V0_3(V0_3),.V0_4(V0_4),.V0_5(V0_5),.V0_6(V0_6),.V0_7(V0_7),
	 .V1_0(V1_0),.V1_1(V1_1),.V1_2(V1_2),.V1_3(V1_3),.V1_4(V1_4),.V1_5(V1_5),.V1_6(V1_6),.V1_7(V1_7),
     .H0_0(H0_0),.H0_1(H0_1),.H0_2(H0_2),.H0_3(H0_3),.H0_4(H0_4),.H0_5(H0_5),.H0_6(H0_6),.H0_7(H0_7),
	 .H1_0(H1_0),.H1_1(H1_1),.H1_2(H1_2),.H1_3(H1_3),.H1_4(H1_4),.H1_5(H1_5),.H1_6(H1_6),.H1_7(H1_7),
      .clk(clk),.reset(reset),.prgm_b(prgm_b),.CLB_prgm_b(CLB_prgm_b),.cb_prgm_b(cb_prgm_b),.sb_prgm_b(sb_prgm_b),.sb_prgm_b_2(sb_prgm_b_2),
	  .bit_in_CLB(bit_in_CLB),.bit_in_CB(bit_in_CB),.sb_prgm_b_in(sb_prgm_b_in),.cb_prgm_b_in(cb_prgm_b_in),.CLB_prgm_b_in(CLB_prgm_b_in),.bit_in_SB(bit_in_SB),.bit_in_SB_2(bit_in_SB_2));


initial begin

CB_config_stream[191:0]= 192'b100000010000001000000100000010000000000000000000_100000010000001000000000000000000010000000000000_000000000000000000000000000000000000000000000000_100000010000001000000100000010000000000000000000;
//CB_config_stream[191:0]= 192'b100000000000000000000000000000000000000000000001_100000000000000000000000000000000000000000000001_100000000000000000000000000000000000000000000001_100000000000000000000000000000000000000000000000;

SB_config_stream[1535:0]= 1536'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_000000000000000011000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
//SB_config_stream[1535:0]= 1536'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001_100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;

SB_config_stream_2[1535:0]= 1536'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

SB_config_stream_3[3071:0]= 3072'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000_000000000000000011000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000011000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

CLB_config_stream[295:0]= 296'b0000000000000000000010000000000000000_0110001101011100000010111111111111111_0000000000000000000010000000000000000_0100001001010100101111000000000000000_0000000000000000000010000000000000000_0000000000000000000010000000000000000_0000000000000000000010000000000000000_0000000001000100001111000000000000000;

for(i=0;i<3072;i=i+1)
SB_config_stream_final[i]=SB_config_stream_3[i];


clk = 1'b0;
 reset=1'b0;
 
 prgm_b=1'b1;   //indicates start of bit_stream----active low
 cb_prgm_b=1'b0;
 sb_prgm_b=1'b0;
  sb_prgm_b_2=1'b0;
 CLB_prgm_b=1'b0;

 fork
 #1 reset=1'b1;
 #1 prgm_b=1'b0;
 #1 cb_prgm_b=1'b1;
  #1 cb_prgm_b_in=1'b1;
   #1 sb_prgm_b=1'b1;
     #1 sb_prgm_b_2=1'b1;
  #1 sb_prgm_b_in=1'b1;
   #1 CLB_prgm_b=1'b1;
  #1 CLB_prgm_b_in=1'b1;

 #1 CB_counter=0;CB_count=0;
  #1 CLB_counter=0;CLB_count=0;
   #1 SB_counter=0;SB_count=0;
      #1 SB_counter_2=0;SB_count_2=0;
 #1 reset=1'b1;
 #2 reset=1'b0;
 join
end



always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && cb_prgm_b!=1'b0) begin

	
	
    if((CB_counter == 49) && cb_prgm_b!=1'b0) //(no of bits required for one CB) + 1= 48+1=49
	begin
	    
		CB_count=CB_count+1;
		
		CB_counter=0;
		if(CB_count==4)
		begin
			
			cb_prgm_b=1'b0;
           // prgm_b=1'b1;
			
		end
	end 
	bit_in_CB <= CB_config_stream[0];
	CB_config_stream <=CB_config_stream>>1;
	CB_counter=CB_counter+1;//if endsj
end 

end //always block ends


always@(posedge clk or posedge reset)
begin 

	if(prgm_b!=1'b1 && sb_prgm_b!=1'b0) begin
	
		if((SB_counter == 769) && sb_prgm_b!=1'b0) //(no of bits required for one SB +1 = 769)
			begin
	    
			SB_count=SB_count+1;
			SB_counter=0;
			if(SB_count==4)
			begin
			
				sb_prgm_b=1'b0;
			sb_prgm_b_in=1'b1;
			 prgm_b=1'b1;
			
			end
		end 
	bit_in_SB <= SB_config_stream_final[0];
	SB_config_stream_final <=SB_config_stream_final>>1;
	SB_counter=SB_counter+1;//if endsj
	end 

end //always block ends
/*
always@(posedge clk or posedge reset)
begin 

	if(prgm_b!=1'b1 && sb_prgm_b_2!=1'b0) begin
	
		if((SB_counter_2 == 769) && sb_prgm_b_2!=1'b0) //(no of bits required for one SB +1 = 769)
			begin
	    
			SB_count_2=SB_count_2+1;
			SB_counter_2=0;
			if(SB_count_2==2)
			begin
			
				sb_prgm_b_2=1'b0;
			sb_prgm_b_in=1'b1;
			if(sb_prgm_b_2==1'b0)
			 	 prgm_b=1'b1;
			
			end
		end 
	bit_in_SB_2 <= SB_config_stream_2[0];
	SB_config_stream_2 <=SB_config_stream_2>>1;
	SB_counter_2=SB_counter_2+1;//if endsj
	end 

end //always block ends  

*/  

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && CLB_prgm_b!=1'b0) 
begin

    if((CLB_counter == 297) && CLB_prgm_b!=1'b0) //(no of bits required for one CLB) + 1= 37+1=38  or (37 + (number of LUT -1))
	begin
	    
		CLB_count=CLB_count+1;
		
		CLB_counter=0;
		if(CLB_count==1)
		begin
			
			CLB_prgm_b=1'b0;
          
			
		end
	end 
	bit_in_CLB <= CLB_config_stream[0];
	CLB_config_stream <=CLB_config_stream>>1;
	CLB_counter=CLB_counter+1;//if endsj
end 

end //always block ends

initial begin
//for(i=0;i<=6074;i++)
//begin

forever #5 clk=!clk;
end

//end

initial
	begin 

	#8350;               //time=5 seconds
V00=1;V01=1;V02=1;V03=1;//H05=1;H06=1;H07=1;H08=1;
H00=0;H01=1;H02=0;H03=1;
//V10=1;V11=1;
#500;
	//reset=1'b0;
V00=1;V01=1;V02=1;V03=1;//H05=1;H06=1;H07=1;H08=1;
H00=0;H01=1;H02=0;H03=1;
//V10=1;V11=1;
	#86500 $finish;
end

initial begin
    $dumpfile("test.vcd");

    $dumpvars(0,FPGA_testbench);
    $timeformat(-9, 1, " ns", 6);
	$monitor("At prgm_b=%b reset=%b SB_count=%d SB_count_2=%d",prgm_b,reset,SB_count,SB_count_2);
end

//Stimulus

endmodule
