
		
	module SB_config_behav(bit_in,prgm_b,clk,reset,sb_prgm_b,N0_E0,N0_E1,N0_E2,N0_E3,N0_E4,N0_E5,N0_E6,N0_E7,N0_S0,N0_S1,N0_S2,N0_S3,N0_S4,N0_S5,N0_S6,N0_S7,N0_W0,N0_W1,N0_W2,N0_W3,N0_W4,N0_W5,N0_W6,N0_W7,N1_E0,
	N1_E1,N1_E2,N1_E3,N1_E4,N1_E5,N1_E6,N1_E7,N1_S0,N1_S1,N1_S2,N1_S3,N1_S4,N1_S5,N1_S6,N1_S7,N1_W0,N1_W1,N1_W2,N1_W3,N1_W4,N1_W5,N1_W6,N1_W7,N2_E0,N2_E1,
	N2_E2,N2_E3,N2_E4,N2_E5,N2_E6,N2_E7,N2_S0,N2_S1,N2_S2,N2_S3,N2_S4,N2_S5,N2_S6,N2_S7,N2_W0,N2_W1,N2_W2,N2_W3,N2_W4,N2_W5,N2_W6,N2_W7,N3_E0,N3_E1,N3_E2,
	N3_E3,N3_E4,N3_E5,N3_E6,N3_E7,N3_S0,N3_S1,N3_S2,N3_S3,N3_S4,N3_S5,N3_S6,N3_S7,N3_W0,N3_W1,N3_W2,N3_W3,N3_W4,N3_W5,N3_W6,N3_W7,N4_E0,N4_E1,N4_E2,N4_E3,
	N4_E4,N4_E5,N4_E6,N4_E7,N4_S0,N4_S1,N4_S2,N4_S3,N4_S4,N4_S5,N4_S6,N4_S7,N4_W0,N4_W1,N4_W2,N4_W3,N4_W4,N4_W5,N4_W6,N4_W7,N5_E0,N5_E1,N5_E2,N5_E3,N5_E4,
	N5_E5,N5_E6,N5_E7,N5_S0,N5_S1,N5_S2,N5_S3,N5_S4,N5_S5,N5_S6,N5_S7,N5_W0,N5_W1,N5_W2,N5_W3,N5_W4,N5_W5,N5_W6,N5_W7,N6_E0,N6_E1,N6_E2,N6_E3,N6_E4,N6_E5,
	N6_E6,N6_E7,N6_S0,N6_S1,N6_S2,N6_S3,N6_S4,N6_S5,N6_S6,N6_S7,N6_W0,N6_W1,N6_W2,N6_W3,N6_W4,N6_W5,N6_W6,N6_W7,N7_E0,N7_E1,N7_E2,N7_E3,N7_E4,N7_E5,N7_E6,
	N7_E7,N7_S0,N7_S1,N7_S2,N7_S3,N7_S4,N7_S5,N7_S6,N7_S7,N7_W0,N7_W1,N7_W2,N7_W3,N7_W4,N7_W5,N7_W6,N7_W7,E0_W0,E0_W1,E0_W2,E0_W3,E0_W4,E0_W5,E0_W6,E0_W7,
	E0_S0,E0_S1,E0_S2,E0_S3,E0_S4,E0_S5,E0_S6,E0_S7,E1_W0,E1_W1,E1_W2,E1_W3,E1_W4,E1_W5,E1_W6,E1_W7,E1_S0,E1_S1,E1_S2,E1_S3,E1_S4,E1_S5,E1_S6,E1_S7,E2_W0,
	E2_W1,E2_W2,E2_W3,E2_W4,E2_W5,E2_W6,E2_W7,E2_S0,E2_S1,E2_S2,E2_S3,E2_S4,E2_S5,E2_S6,E2_S7,E3_W0,E3_W1,E3_W2,E3_W3,E3_W4,E3_W5,E3_W6,E3_W7,E3_S0,E3_S1,
	E3_S2,E3_S3,E3_S4,E3_S5,E3_S6,E3_S7,E4_W0,E4_W1,E4_W2,E4_W3,E4_W4,E4_W5,E4_W6,E4_W7,E4_S0,E4_S1,E4_S2,E4_S3,E4_S4,E4_S5,E4_S6,E4_S7,E5_W0,E5_W1,E5_W2,
	E5_W3,E5_W4,E5_W5,E5_W6,E5_W7,E5_S0,E5_S1,E5_S2,E5_S3,E5_S4,E5_S5,E5_S6,E5_S7,E6_W0,E6_W1,E6_W2,E6_W3,E6_W4,E6_W5,E6_W6,E6_W7,E6_S0,E6_S1,E6_S2,E6_S3,
	E6_S4,E6_S5,E6_S6,E6_S7,E7_W0,E7_W1,E7_W2,E7_W3,E7_W4,E7_W5,E7_W6,E7_W7,E7_S0,E7_S1,E7_S2,E7_S3,E7_S4,E7_S5,E7_S6,E7_S7,S0_W0,S0_W1,S0_W2,S0_W3,S0_W4,
	S0_W5,S0_W6,S0_W7,S1_W0,S1_W1,S1_W2,S1_W3,S1_W4,S1_W5,S1_W6,S1_W7,S2_W0,S2_W1,S2_W2,S2_W3,S2_W4,S2_W5,S2_W6,S2_W7,S3_W0,S3_W1,S3_W2,S3_W3,S3_W4,S3_W5,
	S3_W6,S3_W7,S4_W0,S4_W1,S4_W2,S4_W3,S4_W4,S4_W5,S4_W6,S4_W7,S5_W0,S5_W1,S5_W2,S5_W3,S5_W4,S5_W5,S5_W6,S5_W7,S6_W0,S6_W1,S6_W2,S6_W3,S6_W4,S6_W5,S6_W6,
	S6_W7,S7_W0,S7_W1,S7_W2,S7_W3,S7_W4,S7_W5,S7_W6,S7_W7,sb_prgm_b_in,sb_prgm_b_out);
	input bit_in,prgm_b,sb_prgm_b,sb_prgm_b_in,clk,reset;
	output reg sb_prgm_b_out;
	reg [9:0] count;

	output reg [1:0]N0_E0;output reg [1:0]N0_E1;output reg [1:0]N0_E2;output reg [1:0]N0_E3;output reg [1:0]N0_E4;output reg [1:0]N0_E5;output reg [1:0]N0_E6;output reg [1:0]N0_E7;output reg [1:0]N0_S0;output reg [1:0]N0_S1;output reg [1:0]N0_S2;output reg [1:0]N0_S3;output reg [1:0]N0_S4;output reg [1:0]N0_S5;output reg [1:0]N0_S6;output reg [1:0]N0_S7;output reg [1:0]N0_W0;output reg [1:0]N0_W1;output reg [1:0]N0_W2;output reg [1:0]N0_W3;output reg [1:0]N0_W4;output reg [1:0]N0_W5;output reg [1:0]N0_W6;output reg [1:0]N0_W7;output reg [1:0]N1_E0;
	output reg [1:0]N1_E1;output reg [1:0]N1_E2;output reg [1:0]N1_E3;output reg [1:0]N1_E4;output reg [1:0]N1_E5;output reg [1:0]N1_E6;output reg [1:0]N1_E7;output reg [1:0]N1_S0;output reg [1:0]N1_S1;output reg [1:0]N1_S2;output reg [1:0]N1_S3;output reg [1:0]N1_S4;output reg [1:0]N1_S5;output reg [1:0]N1_S6;output reg [1:0]N1_S7;output reg [1:0]N1_W0;output reg [1:0]N1_W1;output reg [1:0]N1_W2;output reg [1:0]N1_W3;output reg [1:0]N1_W4;output reg [1:0]N1_W5;output reg [1:0]N1_W6;output reg [1:0]N1_W7;output reg [1:0]N2_E0;output reg [1:0]N2_E1;
	output reg [1:0]N2_E2;output reg [1:0]N2_E3;output reg [1:0]N2_E4;output reg [1:0]N2_E5;output reg [1:0]N2_E6;output reg [1:0]N2_E7;output reg [1:0]N2_S0;output reg [1:0]N2_S1;output reg [1:0]N2_S2;output reg [1:0]N2_S3;output reg [1:0]N2_S4;output reg [1:0]N2_S5;output reg [1:0]N2_S6;output reg [1:0]N2_S7;output reg [1:0]N2_W0;output reg [1:0]N2_W1;output reg [1:0]N2_W2;output reg [1:0]N2_W3;output reg [1:0]N2_W4;output reg [1:0]N2_W5;output reg [1:0]N2_W6;output reg [1:0]N2_W7;output reg [1:0]N3_E0;output reg [1:0]N3_E1;output reg [1:0]N3_E2;
	output reg [1:0]N3_E3;output reg [1:0]N3_E4;output reg [1:0]N3_E5;output reg [1:0]N3_E6;output reg [1:0]N3_E7;output reg [1:0]N3_S0;output reg [1:0]N3_S1;output reg [1:0]N3_S2;output reg [1:0]N3_S3;output reg [1:0]N3_S4;output reg [1:0]N3_S5;output reg [1:0]N3_S6;output reg [1:0]N3_S7;output reg [1:0]N3_W0;output reg [1:0]N3_W1;output reg [1:0]N3_W2;output reg [1:0]N3_W3;output reg [1:0]N3_W4;output reg [1:0]N3_W5;output reg [1:0]N3_W6;output reg [1:0]N3_W7;output reg [1:0]N4_E0;output reg [1:0]N4_E1;output reg [1:0]N4_E2;output reg [1:0]N4_E3;
	output reg [1:0]N4_E4;output reg [1:0]N4_E5;output reg [1:0]N4_E6;output reg [1:0]N4_E7;output reg [1:0]N4_S0;output reg [1:0]N4_S1;output reg [1:0]N4_S2;output reg [1:0]N4_S3;output reg [1:0]N4_S4;output reg [1:0]N4_S5;output reg [1:0]N4_S6;output reg [1:0]N4_S7;output reg [1:0]N4_W0;output reg [1:0]N4_W1;output reg [1:0]N4_W2;output reg [1:0]N4_W3;output reg [1:0]N4_W4;output reg [1:0]N4_W5;output reg [1:0]N4_W6;output reg [1:0]N4_W7;output reg [1:0]N5_E0;output reg [1:0]N5_E1;output reg [1:0]N5_E2;output reg [1:0]N5_E3;output reg [1:0]N5_E4;
	output reg [1:0]N5_E5;output reg [1:0]N5_E6;output reg [1:0]N5_E7;output reg [1:0]N5_S0;output reg [1:0]N5_S1;output reg [1:0]N5_S2;output reg [1:0]N5_S3;output reg [1:0]N5_S4;output reg [1:0]N5_S5;output reg [1:0]N5_S6;output reg [1:0]N5_S7;output reg [1:0]N5_W0;output reg [1:0]N5_W1;output reg [1:0]N5_W2;output reg [1:0]N5_W3;output reg [1:0]N5_W4;output reg [1:0]N5_W5;output reg [1:0]N5_W6;output reg [1:0]N5_W7;output reg [1:0]N6_E0;output reg [1:0]N6_E1;output reg [1:0]N6_E2;output reg [1:0]N6_E3;output reg [1:0]N6_E4;output reg [1:0]N6_E5;
	output reg [1:0]N6_E6;output reg [1:0]N6_E7;output reg [1:0]N6_S0;output reg [1:0]N6_S1;output reg [1:0]N6_S2;output reg [1:0]N6_S3;output reg [1:0]N6_S4;output reg [1:0]N6_S5;output reg [1:0]N6_S6;output reg [1:0]N6_S7;output reg [1:0]N6_W0;output reg [1:0]N6_W1;output reg [1:0]N6_W2;output reg [1:0]N6_W3;output reg [1:0]N6_W4;output reg [1:0]N6_W5;output reg [1:0]N6_W6;output reg [1:0]N6_W7;output reg [1:0]N7_E0;output reg [1:0]N7_E1;output reg [1:0]N7_E2;output reg [1:0]N7_E3;output reg [1:0]N7_E4;output reg [1:0]N7_E5;output reg [1:0]N7_E6;
	output reg [1:0]N7_E7;output reg [1:0]N7_S0;output reg [1:0]N7_S1;output reg [1:0]N7_S2;output reg [1:0]N7_S3;output reg [1:0]N7_S4;output reg [1:0]N7_S5;output reg [1:0]N7_S6;output reg [1:0]N7_S7;output reg [1:0]N7_W0;output reg [1:0]N7_W1;output reg [1:0]N7_W2;output reg [1:0]N7_W3;output reg [1:0]N7_W4;output reg [1:0]N7_W5;output reg [1:0]N7_W6;output reg [1:0]N7_W7;output reg [1:0]E0_W0;output reg [1:0]E0_W1;output reg [1:0]E0_W2;output reg [1:0]E0_W3;output reg [1:0]E0_W4;output reg [1:0]E0_W5;output reg [1:0]E0_W6;output reg [1:0]E0_W7;
	output reg [1:0]E0_S0;output reg [1:0]E0_S1;output reg [1:0]E0_S2;output reg [1:0]E0_S3;output reg [1:0]E0_S4;output reg [1:0]E0_S5;output reg [1:0]E0_S6;output reg [1:0]E0_S7;output reg [1:0]E1_W0;output reg [1:0]E1_W1;output reg [1:0]E1_W2;output reg [1:0]E1_W3;output reg [1:0]E1_W4;output reg [1:0]E1_W5;output reg [1:0]E1_W6;output reg [1:0]E1_W7;output reg [1:0]E1_S0;output reg [1:0]E1_S1;output reg [1:0]E1_S2;output reg [1:0]E1_S3;output reg [1:0]E1_S4;output reg [1:0]E1_S5;output reg [1:0]E1_S6;output reg [1:0]E1_S7;output reg [1:0]E2_W0;
	output reg [1:0]E2_W1;output reg [1:0]E2_W2;output reg [1:0]E2_W3;output reg [1:0]E2_W4;output reg [1:0]E2_W5;output reg [1:0]E2_W6;output reg [1:0]E2_W7;output reg [1:0]E2_S0;output reg [1:0]E2_S1;output reg [1:0]E2_S2;output reg [1:0]E2_S3;output reg [1:0]E2_S4;output reg [1:0]E2_S5;output reg [1:0]E2_S6;output reg [1:0]E2_S7;output reg [1:0]E3_W0;output reg [1:0]E3_W1;output reg [1:0]E3_W2;output reg [1:0]E3_W3;output reg [1:0]E3_W4;output reg [1:0]E3_W5;output reg [1:0]E3_W6;output reg [1:0]E3_W7;output reg [1:0]E3_S0;output reg [1:0]E3_S1;
	output reg [1:0]E3_S2;output reg [1:0]E3_S3;output reg [1:0]E3_S4;output reg [1:0]E3_S5;output reg [1:0]E3_S6;output reg [1:0]E3_S7;output reg [1:0]E4_W0;output reg [1:0]E4_W1;output reg [1:0]E4_W2;output reg [1:0]E4_W3;output reg [1:0]E4_W4;output reg [1:0]E4_W5;output reg [1:0]E4_W6;output reg [1:0]E4_W7;output reg [1:0]E4_S0;output reg [1:0]E4_S1;output reg [1:0]E4_S2;output reg [1:0]E4_S3;output reg [1:0]E4_S4;output reg [1:0]E4_S5;output reg [1:0]E4_S6;output reg [1:0]E4_S7;output reg [1:0]E5_W0;output reg [1:0]E5_W1;output reg [1:0]E5_W2;
	output reg [1:0]E5_W3;output reg [1:0]E5_W4;output reg [1:0]E5_W5;output reg [1:0]E5_W6;output reg [1:0]E5_W7;output reg [1:0]E5_S0;output reg [1:0]E5_S1;output reg [1:0]E5_S2;output reg [1:0]E5_S3;output reg [1:0]E5_S4;output reg [1:0]E5_S5;output reg [1:0]E5_S6;output reg [1:0]E5_S7;output reg [1:0]E6_W0;output reg [1:0]E6_W1;output reg [1:0]E6_W2;output reg [1:0]E6_W3;output reg [1:0]E6_W4;output reg [1:0]E6_W5;output reg [1:0]E6_W6;output reg [1:0]E6_W7;output reg [1:0]E6_S0;output reg [1:0]E6_S1;output reg [1:0]E6_S2;output reg [1:0]E6_S3;
	output reg [1:0]E6_S4;output reg [1:0]E6_S5;output reg [1:0]E6_S6;output reg [1:0]E6_S7;output reg [1:0]E7_W0;output reg [1:0]E7_W1;output reg [1:0]E7_W2;output reg [1:0]E7_W3;output reg [1:0]E7_W4;output reg [1:0]E7_W5;output reg [1:0]E7_W6;output reg [1:0]E7_W7;output reg [1:0]E7_S0;output reg [1:0]E7_S1;output reg [1:0]E7_S2;output reg [1:0]E7_S3;output reg [1:0]E7_S4;output reg [1:0]E7_S5;output reg [1:0]E7_S6;output reg [1:0]E7_S7;output reg [1:0]S0_W0;output reg [1:0]S0_W1;output reg [1:0]S0_W2;output reg [1:0]S0_W3;output reg [1:0]S0_W4;
	output reg [1:0]S0_W5;output reg [1:0]S0_W6;output reg [1:0]S0_W7;output reg [1:0]S1_W0;output reg [1:0]S1_W1;output reg [1:0]S1_W2;output reg [1:0]S1_W3;output reg [1:0]S1_W4;output reg [1:0]S1_W5;output reg [1:0]S1_W6;output reg [1:0]S1_W7;output reg [1:0]S2_W0;output reg [1:0]S2_W1;output reg [1:0]S2_W2;output reg [1:0]S2_W3;output reg [1:0]S2_W4;output reg [1:0]S2_W5;output reg [1:0]S2_W6;output reg [1:0]S2_W7;output reg [1:0]S3_W0;output reg [1:0]S3_W1;output reg [1:0]S3_W2;output reg [1:0]S3_W3;output reg [1:0]S3_W4;output reg [1:0]S3_W5;
	output reg [1:0]S3_W6;output reg [1:0]S3_W7;output reg [1:0]S4_W0;output reg [1:0]S4_W1;output reg [1:0]S4_W2;output reg [1:0]S4_W3;output reg [1:0]S4_W4;output reg [1:0]S4_W5;output reg [1:0]S4_W6;output reg [1:0]S4_W7;output reg [1:0]S5_W0;output reg [1:0]S5_W1;output reg [1:0]S5_W2;output reg [1:0]S5_W3;output reg [1:0]S5_W4;output reg [1:0]S5_W5;output reg [1:0]S5_W6;output reg [1:0]S5_W7;output reg [1:0]S6_W0;output reg [1:0]S6_W1;output reg [1:0]S6_W2;output reg [1:0]S6_W3;output reg [1:0]S6_W4;output reg [1:0]S6_W5;output reg [1:0]S6_W6;
	output reg [1:0]S6_W7;output reg [1:0]S7_W0;output reg [1:0]S7_W1;output reg [1:0]S7_W2;output reg [1:0]S7_W3;output reg [1:0]S7_W4;output reg [1:0]S7_W5;output reg [1:0]S7_W6;output reg [1:0]S7_W7;
		
		//output reg bit_out;
	


  initial begin
	count[9:0]=10'b0000000000;
	sb_prgm_b_out=1'b0;
	N0_E0[1:0] <= 2'b00;	 N2_E2[1:0] <= 2'b00;    N4_E4[1:0] <= 2'b00;   N6_E6[1:0] <= 2'b00;   E0_S0[1:0] <= 2'b00;    E3_S2[1:0] <= 2'b00;   E6_S4[1:0] <= 2'b00;   S3_W6[1:0] <= 2'b00;
	N0_E1[1:0] <= 2'b00;     N2_E3[1:0] <= 2'b00;    N4_E5[1:0] <= 2'b00;   N6_E7[1:0] <= 2'b00;   E0_S1[1:0] <= 2'b00;    E3_S3[1:0] <= 2'b00;   E6_S5[1:0] <= 2'b00;   S3_W7[1:0] <= 2'b00;
	N0_E2[1:0] <= 2'b00;     N2_E4[1:0] <= 2'b00;    N4_E6[1:0] <= 2'b00;   N6_S0[1:0] <= 2'b00;   E0_S2[1:0] <= 2'b00;    E3_S4[1:0] <= 2'b00;   E6_S6[1:0] <= 2'b00;   S4_W0[1:0] <= 2'b00;
	N0_E3[1:0] <= 2'b00;     N2_E5[1:0] <= 2'b00;    N4_E7[1:0] <= 2'b00;   N6_S1[1:0] <= 2'b00;   E0_S3[1:0] <= 2'b00;    E3_S5[1:0] <= 2'b00;   E6_S7[1:0] <= 2'b00;   S4_W1[1:0] <= 2'b00;
	N0_E4[1:0] <= 2'b00;     N2_E6[1:0] <= 2'b00;    N4_S0[1:0] <= 2'b00;   N6_S2[1:0] <= 2'b00;   E0_S4[1:0] <= 2'b00;    E3_S6[1:0] <= 2'b00;   E7_W0[1:0] <= 2'b00;   S4_W2[1:0] <= 2'b00;
	N0_E5[1:0] <= 2'b00;     N2_E7[1:0] <= 2'b00;    N4_S1[1:0] <= 2'b00;   N6_S3[1:0] <= 2'b00;   E0_S5[1:0] <= 2'b00;    E3_S7[1:0] <= 2'b00;   E7_W1[1:0] <= 2'b00;   S4_W3[1:0] <= 2'b00;
	N0_E6[1:0] <= 2'b00;     N2_S0[1:0] <= 2'b00;    N4_S2[1:0] <= 2'b00;   N6_S4[1:0] <= 2'b00;   E0_S6[1:0] <= 2'b00;    E4_W0[1:0] <= 2'b00;   E7_W2[1:0] <= 2'b00;   S4_W4[1:0] <= 2'b00;
	N0_E7[1:0] <= 2'b00;     N2_S1[1:0] <= 2'b00;    N4_S3[1:0] <= 2'b00;   N6_S5[1:0] <= 2'b00;   E0_S7[1:0] <= 2'b00;    E4_W1[1:0] <= 2'b00;   E7_W3[1:0] <= 2'b00;   S4_W5[1:0] <= 2'b00;
	N0_S0[1:0] <= 2'b00;     N2_S2[1:0] <= 2'b00;    N4_S4[1:0] <= 2'b00;   N6_S6[1:0] <= 2'b00;   E1_W0[1:0] <= 2'b00;    E4_W2[1:0] <= 2'b00;   E7_W4[1:0] <= 2'b00;   S4_W6[1:0] <= 2'b00;
	N0_S1[1:0] <= 2'b00;     N2_S3[1:0] <= 2'b00;    N4_S5[1:0] <= 2'b00;   N6_S7[1:0] <= 2'b00;   E1_W1[1:0] <= 2'b00;    E4_W3[1:0] <= 2'b00;   E7_W5[1:0] <= 2'b00;   S4_W7[1:0] <= 2'b00;
	N0_S2[1:0] <= 2'b00;     N2_S4[1:0] <= 2'b00;    N4_S6[1:0] <= 2'b00;   N6_W0[1:0] <= 2'b00;   E1_W2[1:0] <= 2'b00;    E4_W4[1:0] <= 2'b00;   E7_W6[1:0] <= 2'b00;   S5_W0[1:0] <= 2'b00;
	N0_S3[1:0] <= 2'b00;     N2_S5[1:0] <= 2'b00;    N4_S7[1:0] <= 2'b00;   N6_W1[1:0] <= 2'b00;   E1_W3[1:0] <= 2'b00;    E4_W5[1:0] <= 2'b00;   E7_W7[1:0] <= 2'b00;   S5_W1[1:0] <= 2'b00;
	N0_S4[1:0] <= 2'b00;     N2_S6[1:0] <= 2'b00;    N4_W0[1:0] <= 2'b00;   N6_W2[1:0] <= 2'b00;   E1_W4[1:0] <= 2'b00;    E4_W6[1:0] <= 2'b00;   E7_S0[1:0] <= 2'b00;   S5_W2[1:0] <= 2'b00;
	N0_S5[1:0] <= 2'b00;     N2_S7[1:0] <= 2'b00;    N4_W1[1:0] <= 2'b00;   N6_W3[1:0] <= 2'b00;   E1_W5[1:0] <= 2'b00;    E4_W7[1:0] <= 2'b00;   E7_S1[1:0] <= 2'b00;   S5_W3[1:0] <= 2'b00;
	N0_S6[1:0] <= 2'b00;     N2_W0[1:0] <= 2'b00;    N4_W2[1:0] <= 2'b00;   N6_W4[1:0] <= 2'b00;   E1_W6[1:0] <= 2'b00;    E4_S0[1:0] <= 2'b00;   E7_S2[1:0] <= 2'b00;   S5_W4[1:0] <= 2'b00;
	N0_S7[1:0] <= 2'b00;     N2_W1[1:0] <= 2'b00;    N4_W3[1:0] <= 2'b00;   N6_W5[1:0] <= 2'b00;   E1_W7[1:0] <= 2'b00;    E4_S1[1:0] <= 2'b00;   E7_S3[1:0] <= 2'b00;   S5_W5[1:0] <= 2'b00;
	N0_W0[1:0] <= 2'b00;     N2_W2[1:0] <= 2'b00;    N4_W4[1:0] <= 2'b00;   N6_W6[1:0] <= 2'b00;   E1_S0[1:0] <= 2'b00;    E4_S2[1:0] <= 2'b00;   E7_S4[1:0] <= 2'b00;   S5_W6[1:0] <= 2'b00;
	N0_W1[1:0] <= 2'b00;     N2_W3[1:0] <= 2'b00;    N4_W5[1:0] <= 2'b00;   N6_W7[1:0] <= 2'b00;   E1_S1[1:0] <= 2'b00;    E4_S3[1:0] <= 2'b00;   E7_S5[1:0] <= 2'b00;   S5_W7[1:0] <= 2'b00;
	N0_W2[1:0] <= 2'b00;     N2_W4[1:0] <= 2'b00;    N4_W6[1:0] <= 2'b00;   N7_E0[1:0] <= 2'b00;   E1_S2[1:0] <= 2'b00;    E4_S4[1:0] <= 2'b00;   E7_S6[1:0] <= 2'b00;   S6_W0[1:0] <= 2'b00;
	N0_W3[1:0] <= 2'b00;     N2_W5[1:0] <= 2'b00;    N4_W7[1:0] <= 2'b00;   N7_E1[1:0] <= 2'b00;   E1_S3[1:0] <= 2'b00;    E4_S5[1:0] <= 2'b00;   E7_S7[1:0] <= 2'b00;   S6_W1[1:0] <= 2'b00;
	N0_W4[1:0] <= 2'b00;     N2_W6[1:0] <= 2'b00;    N5_E0[1:0] <= 2'b00;   N7_E2[1:0] <= 2'b00;   E1_S4[1:0] <= 2'b00;    E4_S6[1:0] <= 2'b00;   S0_W0[1:0] <= 2'b00;   S6_W2[1:0] <= 2'b00;
	N0_W5[1:0] <= 2'b00;     N2_W7[1:0] <= 2'b00;    N5_E1[1:0] <= 2'b00;   N7_E3[1:0] <= 2'b00;   E1_S5[1:0] <= 2'b00;    E4_S7[1:0] <= 2'b00;   S0_W1[1:0] <= 2'b00;   S6_W3[1:0] <= 2'b00;
	N0_W6[1:0] <= 2'b00;     N3_E0[1:0] <= 2'b00;    N5_E2[1:0] <= 2'b00;   N7_E4[1:0] <= 2'b00;   E1_S6[1:0] <= 2'b00;    E5_W0[1:0] <= 2'b00;   S0_W2[1:0] <= 2'b00;   S6_W4[1:0] <= 2'b00;
	N0_W7[1:0] <= 2'b00;     N3_E1[1:0] <= 2'b00;    N5_E3[1:0] <= 2'b00;   N7_E5[1:0] <= 2'b00;   E1_S7[1:0] <= 2'b00;    E5_W1[1:0] <= 2'b00;   S0_W3[1:0] <= 2'b00;   S6_W5[1:0] <= 2'b00;
	N1_E0[1:0] <= 2'b00;     N3_E2[1:0] <= 2'b00;    N5_E4[1:0] <= 2'b00;   N7_E6[1:0] <= 2'b00;   E2_W0[1:0] <= 2'b00;    E5_W2[1:0] <= 2'b00;   S0_W4[1:0] <= 2'b00;   S6_W6[1:0] <= 2'b00;
	N1_E1[1:0] <= 2'b00;     N3_E3[1:0] <= 2'b00;    N5_E5[1:0] <= 2'b00;   N7_E7[1:0] <= 2'b00;   E2_W1[1:0] <= 2'b00;    E5_W3[1:0] <= 2'b00;   S0_W5[1:0] <= 2'b00;   S6_W7[1:0] <= 2'b00;
	N1_E2[1:0] <= 2'b00;     N3_E4[1:0] <= 2'b00;    N5_E6[1:0] <= 2'b00;   N7_S0[1:0] <= 2'b00;   E2_W2[1:0] <= 2'b00;    E5_W4[1:0] <= 2'b00;   S0_W6[1:0] <= 2'b00;   S7_W0[1:0] <= 2'b00;
	N1_E3[1:0] <= 2'b00;     N3_E5[1:0] <= 2'b00;    N5_E7[1:0] <= 2'b00;   N7_S1[1:0] <= 2'b00;   E2_W3[1:0] <= 2'b00;    E5_W5[1:0] <= 2'b00;   S0_W7[1:0] <= 2'b00;   S7_W1[1:0] <= 2'b00;
	N1_E4[1:0] <= 2'b00;     N3_E6[1:0] <= 2'b00;    N5_S0[1:0] <= 2'b00;   N7_S2[1:0] <= 2'b00;   E2_W4[1:0] <= 2'b00;    E5_W6[1:0] <= 2'b00;   S1_W0[1:0] <= 2'b00;   S7_W2[1:0] <= 2'b00;
	N1_E5[1:0] <= 2'b00;     N3_E7[1:0] <= 2'b00;    N5_S1[1:0] <= 2'b00;   N7_S3[1:0] <= 2'b00;   E2_W5[1:0] <= 2'b00;    E5_W7[1:0] <= 2'b00;   S1_W1[1:0] <= 2'b00;   S7_W3[1:0] <= 2'b00;
	N1_E6[1:0] <= 2'b00;     N3_S0[1:0] <= 2'b00;    N5_S2[1:0] <= 2'b00;   N7_S4[1:0] <= 2'b00;   E2_W6[1:0] <= 2'b00;    E5_S0[1:0] <= 2'b00;   S1_W2[1:0] <= 2'b00;   S7_W4[1:0] <= 2'b00;
	N1_E7[1:0] <= 2'b00;     N3_S1[1:0] <= 2'b00;    N5_S3[1:0] <= 2'b00;   N7_S5[1:0] <= 2'b00;   E2_W7[1:0] <= 2'b00;    E5_S1[1:0] <= 2'b00;   S1_W3[1:0] <= 2'b00;   S7_W5[1:0] <= 2'b00;
	N1_S0[1:0] <= 2'b00;     N3_S2[1:0] <= 2'b00;    N5_S4[1:0] <= 2'b00;   N7_S6[1:0] <= 2'b00;   E2_S0[1:0] <= 2'b00;    E5_S2[1:0] <= 2'b00;   S1_W4[1:0] <= 2'b00;   S7_W6[1:0] <= 2'b00;
	N1_S1[1:0] <= 2'b00;     N3_S3[1:0] <= 2'b00;    N5_S5[1:0] <= 2'b00;   N7_S7[1:0] <= 2'b00;   E2_S1[1:0] <= 2'b00;    E5_S3[1:0] <= 2'b00;   S1_W5[1:0] <= 2'b00;   S7_W7[1:0] <= 2'b00;
	N1_S2[1:0] <= 2'b00;     N3_S4[1:0] <= 2'b00;    N5_S6[1:0] <= 2'b00;   N7_W0[1:0] <= 2'b00;   E2_S2[1:0] <= 2'b00;    E5_S4[1:0] <= 2'b00;   S1_W6[1:0] <= 2'b00;  
	N1_S3[1:0] <= 2'b00;     N3_S5[1:0] <= 2'b00;    N5_S7[1:0] <= 2'b00;   N7_W1[1:0] <= 2'b00;   E2_S3[1:0] <= 2'b00;    E5_S5[1:0] <= 2'b00;   S1_W7[1:0] <= 2'b00;
	N1_S4[1:0] <= 2'b00;     N3_S6[1:0] <= 2'b00;    N5_W0[1:0] <= 2'b00;   N7_W2[1:0] <= 2'b00;   E2_S4[1:0] <= 2'b00;    E5_S6[1:0] <= 2'b00;   S2_W0[1:0] <= 2'b00;
	N1_S5[1:0] <= 2'b00;     N3_S7[1:0] <= 2'b00;    N5_W1[1:0] <= 2'b00;   N7_W3[1:0] <= 2'b00;   E2_S5[1:0] <= 2'b00;    E5_S7[1:0] <= 2'b00;   S2_W1[1:0] <= 2'b00;
	N1_S6[1:0] <= 2'b00;     N3_W0[1:0] <= 2'b00;    N5_W2[1:0] <= 2'b00;   N7_W4[1:0] <= 2'b00;   E2_S6[1:0] <= 2'b00;    E6_W0[1:0] <= 2'b00;   S2_W2[1:0] <= 2'b00;
	N1_S7[1:0] <= 2'b00;     N3_W1[1:0] <= 2'b00;    N5_W3[1:0] <= 2'b00;   N7_W5[1:0] <= 2'b00;   E2_S7[1:0] <= 2'b00;    E6_W1[1:0] <= 2'b00;   S2_W3[1:0] <= 2'b00;
	N1_W0[1:0] <= 2'b00;     N3_W2[1:0] <= 2'b00;    N5_W4[1:0] <= 2'b00;   N7_W6[1:0] <= 2'b00;   E3_W0[1:0] <= 2'b00;    E6_W2[1:0] <= 2'b00;   S2_W4[1:0] <= 2'b00;
	N1_W1[1:0] <= 2'b00;     N3_W3[1:0] <= 2'b00;    N5_W5[1:0] <= 2'b00;   N7_W7[1:0] <= 2'b00;   E3_W1[1:0] <= 2'b00;    E6_W3[1:0] <= 2'b00;   S2_W5[1:0] <= 2'b00;
	N1_W2[1:0] <= 2'b00;     N3_W4[1:0] <= 2'b00;    N5_W6[1:0] <= 2'b00;   E0_W0[1:0] <= 2'b00;   E3_W2[1:0] <= 2'b00;    E6_W4[1:0] <= 2'b00;   S2_W6[1:0] <= 2'b00;
	N1_W3[1:0] <= 2'b00;     N3_W5[1:0] <= 2'b00;    N5_W7[1:0] <= 2'b00;   E0_W1[1:0] <= 2'b00;   E3_W3[1:0] <= 2'b00;    E6_W5[1:0] <= 2'b00;   S2_W7[1:0] <= 2'b00;
	N1_W4[1:0] <= 2'b00;     N3_W6[1:0] <= 2'b00;    N6_E0[1:0] <= 2'b00;   E0_W2[1:0] <= 2'b00;   E3_W4[1:0] <= 2'b00;    E6_W6[1:0] <= 2'b00;   S3_W0[1:0] <= 2'b00;
	N1_W5[1:0] <= 2'b00;     N3_W7[1:0] <= 2'b00;    N6_E1[1:0] <= 2'b00;   E0_W3[1:0] <= 2'b00;   E3_W5[1:0] <= 2'b00;    E6_W7[1:0] <= 2'b00;   S3_W1[1:0] <= 2'b00;
	N1_W6[1:0] <= 2'b00;     N4_E0[1:0] <= 2'b00;    N6_E2[1:0] <= 2'b00;   E0_W4[1:0] <= 2'b00;   E3_W6[1:0] <= 2'b00;    E6_S0[1:0] <= 2'b00;   S3_W2[1:0] <= 2'b00;
	N1_W7[1:0] <= 2'b00;     N4_E1[1:0] <= 2'b00;    N6_E3[1:0] <= 2'b00;   E0_W5[1:0] <= 2'b00;   E3_W7[1:0] <= 2'b00;    E6_S1[1:0] <= 2'b00;   S3_W3[1:0] <= 2'b00;
	N2_E0[1:0] <= 2'b00;     N4_E2[1:0] <= 2'b00;    N6_E4[1:0] <= 2'b00;   E0_W6[1:0] <= 2'b00;   E3_S0[1:0] <= 2'b00;    E6_S2[1:0] <= 2'b00;   S3_W4[1:0] <= 2'b00;
	N2_E1[1:0] <= 2'b00;     N4_E3[1:0] <= 2'b00;    N6_E5[1:0] <= 2'b00;   E0_W7[1:0] <= 2'b00;   E3_S1[1:0] <= 2'b00;    E6_S3[1:0] <= 2'b00;   S3_W5[1:0] <= 2'b00;

end

always @(posedge clk or posedge reset)
 begin
	if(prgm_b==1'b0 && sb_prgm_b_in==1'b1 && sb_prgm_b_out!=1'b1 && sb_prgm_b==1'b1)	
	begin
	if(reset)
		sb_prgm_b_out=1'b0;
		
	else begin
		count[9:0]=count[9:0]+1'b1; 
		if(count[9:0]==10'b1100000000)
		begin
			sb_prgm_b_out= 1'b1;
			count[9:0]=10'b0000000000;
			//prgm_b_out=1'b0;
		end  //ends
	end //else ends

	
	end	 //first if ends

end //always block ends




	always @ (posedge clk or posedge reset)
	begin
	if (prgm_b==1'b0 && sb_prgm_b_in==1'b1 && sb_prgm_b_out!=1'b1 && sb_prgm_b==1'b1) begin
	if(reset) begin
	N0_E0[1:0] <= 2'b00;	 N2_E2[1:0] <= 2'b00;    N4_E4[1:0] <= 2'b00;   N6_E6[1:0] <= 2'b00;   E0_S0[1:0] <= 2'b00;    E3_S2[1:0] <= 2'b00;   E6_S4[1:0] <= 2'b00;   S3_W6[1:0] <= 2'b00;
	N0_E1[1:0] <= 2'b00;     N2_E3[1:0] <= 2'b00;    N4_E5[1:0] <= 2'b00;   N6_E7[1:0] <= 2'b00;   E0_S1[1:0] <= 2'b00;    E3_S3[1:0] <= 2'b00;   E6_S5[1:0] <= 2'b00;   S3_W7[1:0] <= 2'b00;
	N0_E2[1:0] <= 2'b00;     N2_E4[1:0] <= 2'b00;    N4_E6[1:0] <= 2'b00;   N6_S0[1:0] <= 2'b00;   E0_S2[1:0] <= 2'b00;    E3_S4[1:0] <= 2'b00;   E6_S6[1:0] <= 2'b00;   S4_W0[1:0] <= 2'b00;
	N0_E3[1:0] <= 2'b00;     N2_E5[1:0] <= 2'b00;    N4_E7[1:0] <= 2'b00;   N6_S1[1:0] <= 2'b00;   E0_S3[1:0] <= 2'b00;    E3_S5[1:0] <= 2'b00;   E6_S7[1:0] <= 2'b00;   S4_W1[1:0] <= 2'b00;
	N0_E4[1:0] <= 2'b00;     N2_E6[1:0] <= 2'b00;    N4_S0[1:0] <= 2'b00;   N6_S2[1:0] <= 2'b00;   E0_S4[1:0] <= 2'b00;    E3_S6[1:0] <= 2'b00;   E7_W0[1:0] <= 2'b00;   S4_W2[1:0] <= 2'b00;
	N0_E5[1:0] <= 2'b00;     N2_E7[1:0] <= 2'b00;    N4_S1[1:0] <= 2'b00;   N6_S3[1:0] <= 2'b00;   E0_S5[1:0] <= 2'b00;    E3_S7[1:0] <= 2'b00;   E7_W1[1:0] <= 2'b00;   S4_W3[1:0] <= 2'b00;
	N0_E6[1:0] <= 2'b00;     N2_S0[1:0] <= 2'b00;    N4_S2[1:0] <= 2'b00;   N6_S4[1:0] <= 2'b00;   E0_S6[1:0] <= 2'b00;    E4_W0[1:0] <= 2'b00;   E7_W2[1:0] <= 2'b00;   S4_W4[1:0] <= 2'b00;
	N0_E7[1:0] <= 2'b00;     N2_S1[1:0] <= 2'b00;    N4_S3[1:0] <= 2'b00;   N6_S5[1:0] <= 2'b00;   E0_S7[1:0] <= 2'b00;    E4_W1[1:0] <= 2'b00;   E7_W3[1:0] <= 2'b00;   S4_W5[1:0] <= 2'b00;
	N0_S0[1:0] <= 2'b00;     N2_S2[1:0] <= 2'b00;    N4_S4[1:0] <= 2'b00;   N6_S6[1:0] <= 2'b00;   E1_W0[1:0] <= 2'b00;    E4_W2[1:0] <= 2'b00;   E7_W4[1:0] <= 2'b00;   S4_W6[1:0] <= 2'b00;
	N0_S1[1:0] <= 2'b00;     N2_S3[1:0] <= 2'b00;    N4_S5[1:0] <= 2'b00;   N6_S7[1:0] <= 2'b00;   E1_W1[1:0] <= 2'b00;    E4_W3[1:0] <= 2'b00;   E7_W5[1:0] <= 2'b00;   S4_W7[1:0] <= 2'b00;
	N0_S2[1:0] <= 2'b00;     N2_S4[1:0] <= 2'b00;    N4_S6[1:0] <= 2'b00;   N6_W0[1:0] <= 2'b00;   E1_W2[1:0] <= 2'b00;    E4_W4[1:0] <= 2'b00;   E7_W6[1:0] <= 2'b00;   S5_W0[1:0] <= 2'b00;
	N0_S3[1:0] <= 2'b00;     N2_S5[1:0] <= 2'b00;    N4_S7[1:0] <= 2'b00;   N6_W1[1:0] <= 2'b00;   E1_W3[1:0] <= 2'b00;    E4_W5[1:0] <= 2'b00;   E7_W7[1:0] <= 2'b00;   S5_W1[1:0] <= 2'b00;
	N0_S4[1:0] <= 2'b00;     N2_S6[1:0] <= 2'b00;    N4_W0[1:0] <= 2'b00;   N6_W2[1:0] <= 2'b00;   E1_W4[1:0] <= 2'b00;    E4_W6[1:0] <= 2'b00;   E7_S0[1:0] <= 2'b00;   S5_W2[1:0] <= 2'b00;
	N0_S5[1:0] <= 2'b00;     N2_S7[1:0] <= 2'b00;    N4_W1[1:0] <= 2'b00;   N6_W3[1:0] <= 2'b00;   E1_W5[1:0] <= 2'b00;    E4_W7[1:0] <= 2'b00;   E7_S1[1:0] <= 2'b00;   S5_W3[1:0] <= 2'b00;
	N0_S6[1:0] <= 2'b00;     N2_W0[1:0] <= 2'b00;    N4_W2[1:0] <= 2'b00;   N6_W4[1:0] <= 2'b00;   E1_W6[1:0] <= 2'b00;    E4_S0[1:0] <= 2'b00;   E7_S2[1:0] <= 2'b00;   S5_W4[1:0] <= 2'b00;
	N0_S7[1:0] <= 2'b00;     N2_W1[1:0] <= 2'b00;    N4_W3[1:0] <= 2'b00;   N6_W5[1:0] <= 2'b00;   E1_W7[1:0] <= 2'b00;    E4_S1[1:0] <= 2'b00;   E7_S3[1:0] <= 2'b00;   S5_W5[1:0] <= 2'b00;
	N0_W0[1:0] <= 2'b00;     N2_W2[1:0] <= 2'b00;    N4_W4[1:0] <= 2'b00;   N6_W6[1:0] <= 2'b00;   E1_S0[1:0] <= 2'b00;    E4_S2[1:0] <= 2'b00;   E7_S4[1:0] <= 2'b00;   S5_W6[1:0] <= 2'b00;
	N0_W1[1:0] <= 2'b00;     N2_W3[1:0] <= 2'b00;    N4_W5[1:0] <= 2'b00;   N6_W7[1:0] <= 2'b00;   E1_S1[1:0] <= 2'b00;    E4_S3[1:0] <= 2'b00;   E7_S5[1:0] <= 2'b00;   S5_W7[1:0] <= 2'b00;
	N0_W2[1:0] <= 2'b00;     N2_W4[1:0] <= 2'b00;    N4_W6[1:0] <= 2'b00;   N7_E0[1:0] <= 2'b00;   E1_S2[1:0] <= 2'b00;    E4_S4[1:0] <= 2'b00;   E7_S6[1:0] <= 2'b00;   S6_W0[1:0] <= 2'b00;
	N0_W3[1:0] <= 2'b00;     N2_W5[1:0] <= 2'b00;    N4_W7[1:0] <= 2'b00;   N7_E1[1:0] <= 2'b00;   E1_S3[1:0] <= 2'b00;    E4_S5[1:0] <= 2'b00;   E7_S7[1:0] <= 2'b00;   S6_W1[1:0] <= 2'b00;
	N0_W4[1:0] <= 2'b00;     N2_W6[1:0] <= 2'b00;    N5_E0[1:0] <= 2'b00;   N7_E2[1:0] <= 2'b00;   E1_S4[1:0] <= 2'b00;    E4_S6[1:0] <= 2'b00;   S0_W0[1:0] <= 2'b00;   S6_W2[1:0] <= 2'b00;
	N0_W5[1:0] <= 2'b00;     N2_W7[1:0] <= 2'b00;    N5_E1[1:0] <= 2'b00;   N7_E3[1:0] <= 2'b00;   E1_S5[1:0] <= 2'b00;    E4_S7[1:0] <= 2'b00;   S0_W1[1:0] <= 2'b00;   S6_W3[1:0] <= 2'b00;
	N0_W6[1:0] <= 2'b00;     N3_E0[1:0] <= 2'b00;    N5_E2[1:0] <= 2'b00;   N7_E4[1:0] <= 2'b00;   E1_S6[1:0] <= 2'b00;    E5_W0[1:0] <= 2'b00;   S0_W2[1:0] <= 2'b00;   S6_W4[1:0] <= 2'b00;
	N0_W7[1:0] <= 2'b00;     N3_E1[1:0] <= 2'b00;    N5_E3[1:0] <= 2'b00;   N7_E5[1:0] <= 2'b00;   E1_S7[1:0] <= 2'b00;    E5_W1[1:0] <= 2'b00;   S0_W3[1:0] <= 2'b00;   S6_W5[1:0] <= 2'b00;
	N1_E0[1:0] <= 2'b00;     N3_E2[1:0] <= 2'b00;    N5_E4[1:0] <= 2'b00;   N7_E6[1:0] <= 2'b00;   E2_W0[1:0] <= 2'b00;    E5_W2[1:0] <= 2'b00;   S0_W4[1:0] <= 2'b00;   S6_W6[1:0] <= 2'b00;
	N1_E1[1:0] <= 2'b00;     N3_E3[1:0] <= 2'b00;    N5_E5[1:0] <= 2'b00;   N7_E7[1:0] <= 2'b00;   E2_W1[1:0] <= 2'b00;    E5_W3[1:0] <= 2'b00;   S0_W5[1:0] <= 2'b00;   S6_W7[1:0] <= 2'b00;
	N1_E2[1:0] <= 2'b00;     N3_E4[1:0] <= 2'b00;    N5_E6[1:0] <= 2'b00;   N7_S0[1:0] <= 2'b00;   E2_W2[1:0] <= 2'b00;    E5_W4[1:0] <= 2'b00;   S0_W6[1:0] <= 2'b00;   S7_W0[1:0] <= 2'b00;
	N1_E3[1:0] <= 2'b00;     N3_E5[1:0] <= 2'b00;    N5_E7[1:0] <= 2'b00;   N7_S1[1:0] <= 2'b00;   E2_W3[1:0] <= 2'b00;    E5_W5[1:0] <= 2'b00;   S0_W7[1:0] <= 2'b00;   S7_W1[1:0] <= 2'b00;
	N1_E4[1:0] <= 2'b00;     N3_E6[1:0] <= 2'b00;    N5_S0[1:0] <= 2'b00;   N7_S2[1:0] <= 2'b00;   E2_W4[1:0] <= 2'b00;    E5_W6[1:0] <= 2'b00;   S1_W0[1:0] <= 2'b00;   S7_W2[1:0] <= 2'b00;
	N1_E5[1:0] <= 2'b00;     N3_E7[1:0] <= 2'b00;    N5_S1[1:0] <= 2'b00;   N7_S3[1:0] <= 2'b00;   E2_W5[1:0] <= 2'b00;    E5_W7[1:0] <= 2'b00;   S1_W1[1:0] <= 2'b00;   S7_W3[1:0] <= 2'b00;
	N1_E6[1:0] <= 2'b00;     N3_S0[1:0] <= 2'b00;    N5_S2[1:0] <= 2'b00;   N7_S4[1:0] <= 2'b00;   E2_W6[1:0] <= 2'b00;    E5_S0[1:0] <= 2'b00;   S1_W2[1:0] <= 2'b00;   S7_W4[1:0] <= 2'b00;
	N1_E7[1:0] <= 2'b00;     N3_S1[1:0] <= 2'b00;    N5_S3[1:0] <= 2'b00;   N7_S5[1:0] <= 2'b00;   E2_W7[1:0] <= 2'b00;    E5_S1[1:0] <= 2'b00;   S1_W3[1:0] <= 2'b00;   S7_W5[1:0] <= 2'b00;
	N1_S0[1:0] <= 2'b00;     N3_S2[1:0] <= 2'b00;    N5_S4[1:0] <= 2'b00;   N7_S6[1:0] <= 2'b00;   E2_S0[1:0] <= 2'b00;    E5_S2[1:0] <= 2'b00;   S1_W4[1:0] <= 2'b00;   S7_W6[1:0] <= 2'b00;
	N1_S1[1:0] <= 2'b00;     N3_S3[1:0] <= 2'b00;    N5_S5[1:0] <= 2'b00;   N7_S7[1:0] <= 2'b00;   E2_S1[1:0] <= 2'b00;    E5_S3[1:0] <= 2'b00;   S1_W5[1:0] <= 2'b00;   S7_W7[1:0] <= 2'b00;
	N1_S2[1:0] <= 2'b00;     N3_S4[1:0] <= 2'b00;    N5_S6[1:0] <= 2'b00;   N7_W0[1:0] <= 2'b00;   E2_S2[1:0] <= 2'b00;    E5_S4[1:0] <= 2'b00;   S1_W6[1:0] <= 2'b00;  
	N1_S3[1:0] <= 2'b00;     N3_S5[1:0] <= 2'b00;    N5_S7[1:0] <= 2'b00;   N7_W1[1:0] <= 2'b00;   E2_S3[1:0] <= 2'b00;    E5_S5[1:0] <= 2'b00;   S1_W7[1:0] <= 2'b00;
	N1_S4[1:0] <= 2'b00;     N3_S6[1:0] <= 2'b00;    N5_W0[1:0] <= 2'b00;   N7_W2[1:0] <= 2'b00;   E2_S4[1:0] <= 2'b00;    E5_S6[1:0] <= 2'b00;   S2_W0[1:0] <= 2'b00;
	N1_S5[1:0] <= 2'b00;     N3_S7[1:0] <= 2'b00;    N5_W1[1:0] <= 2'b00;   N7_W3[1:0] <= 2'b00;   E2_S5[1:0] <= 2'b00;    E5_S7[1:0] <= 2'b00;   S2_W1[1:0] <= 2'b00;
	N1_S6[1:0] <= 2'b00;     N3_W0[1:0] <= 2'b00;    N5_W2[1:0] <= 2'b00;   N7_W4[1:0] <= 2'b00;   E2_S6[1:0] <= 2'b00;    E6_W0[1:0] <= 2'b00;   S2_W2[1:0] <= 2'b00;
	N1_S7[1:0] <= 2'b00;     N3_W1[1:0] <= 2'b00;    N5_W3[1:0] <= 2'b00;   N7_W5[1:0] <= 2'b00;   E2_S7[1:0] <= 2'b00;    E6_W1[1:0] <= 2'b00;   S2_W3[1:0] <= 2'b00;
	N1_W0[1:0] <= 2'b00;     N3_W2[1:0] <= 2'b00;    N5_W4[1:0] <= 2'b00;   N7_W6[1:0] <= 2'b00;   E3_W0[1:0] <= 2'b00;    E6_W2[1:0] <= 2'b00;   S2_W4[1:0] <= 2'b00;
	N1_W1[1:0] <= 2'b00;     N3_W3[1:0] <= 2'b00;    N5_W5[1:0] <= 2'b00;   N7_W7[1:0] <= 2'b00;   E3_W1[1:0] <= 2'b00;    E6_W3[1:0] <= 2'b00;   S2_W5[1:0] <= 2'b00;
	N1_W2[1:0] <= 2'b00;     N3_W4[1:0] <= 2'b00;    N5_W6[1:0] <= 2'b00;   E0_W0[1:0] <= 2'b00;   E3_W2[1:0] <= 2'b00;    E6_W4[1:0] <= 2'b00;   S2_W6[1:0] <= 2'b00;
	N1_W3[1:0] <= 2'b00;     N3_W5[1:0] <= 2'b00;    N5_W7[1:0] <= 2'b00;   E0_W1[1:0] <= 2'b00;   E3_W3[1:0] <= 2'b00;    E6_W5[1:0] <= 2'b00;   S2_W7[1:0] <= 2'b00;
	N1_W4[1:0] <= 2'b00;     N3_W6[1:0] <= 2'b00;    N6_E0[1:0] <= 2'b00;   E0_W2[1:0] <= 2'b00;   E3_W4[1:0] <= 2'b00;    E6_W6[1:0] <= 2'b00;   S3_W0[1:0] <= 2'b00;
	N1_W5[1:0] <= 2'b00;     N3_W7[1:0] <= 2'b00;    N6_E1[1:0] <= 2'b00;   E0_W3[1:0] <= 2'b00;   E3_W5[1:0] <= 2'b00;    E6_W7[1:0] <= 2'b00;   S3_W1[1:0] <= 2'b00;
	N1_W6[1:0] <= 2'b00;     N4_E0[1:0] <= 2'b00;    N6_E2[1:0] <= 2'b00;   E0_W4[1:0] <= 2'b00;   E3_W6[1:0] <= 2'b00;    E6_S0[1:0] <= 2'b00;   S3_W2[1:0] <= 2'b00;
	N1_W7[1:0] <= 2'b00;     N4_E1[1:0] <= 2'b00;    N6_E3[1:0] <= 2'b00;   E0_W5[1:0] <= 2'b00;   E3_W7[1:0] <= 2'b00;    E6_S1[1:0] <= 2'b00;   S3_W3[1:0] <= 2'b00;
	N2_E0[1:0] <= 2'b00;     N4_E2[1:0] <= 2'b00;    N6_E4[1:0] <= 2'b00;   E0_W6[1:0] <= 2'b00;   E3_S0[1:0] <= 2'b00;    E6_S2[1:0] <= 2'b00;   S3_W4[1:0] <= 2'b00;
	N2_E1[1:0] <= 2'b00;     N4_E3[1:0] <= 2'b00;    N6_E5[1:0] <= 2'b00;   E0_W7[1:0] <= 2'b00;   E3_S1[1:0] <= 2'b00;    E6_S3[1:0] <= 2'b00;   S3_W5[1:0] <= 2'b00;

  

	end
	else begin
	N0_E0[1] <= bit_in  ;    N2_E2[1] <= N2_E1[0];   N4_E4[1] <= N4_E3[0];   N6_E6[1] <= N6_E5[0];   E0_S0[1] <= E0_W7[0];   E3_S2[1] <= E3_S1[0];   E6_S4[1] <= E6_S3[0]; S3_W6[1] <= S3_W5[0];
	N0_E0[0] <= N0_E0[1];    N2_E2[0] <= N2_E2[1];   N4_E4[0] <= N4_E4[1];   N6_E6[0] <= N6_E6[1];   E0_S0[0] <= E0_S0[1];   E3_S2[0] <= E3_S2[1];   E6_S4[0] <= E6_S4[1]; S3_W6[0] <= S3_W6[1];
	N0_E1[1] <= N0_E0[0];    N2_E3[1] <= N2_E2[0];   N4_E5[1] <= N4_E4[0];   N6_E7[1] <= N6_E6[0];   E0_S1[1] <= E0_S0[0];   E3_S3[1] <= E3_S2[0];   E6_S5[1] <= E6_S4[0]; S3_W7[1] <= S3_W6[0];
	N0_E1[0] <= N0_E1[1];    N2_E3[0] <= N2_E3[1];   N4_E5[0] <= N4_E5[1];   N6_E7[0] <= N6_E7[1];   E0_S1[0] <= E0_S1[1];   E3_S3[0] <= E3_S3[1];   E6_S5[0] <= E6_S5[1]; S3_W7[0] <= S3_W7[1];
	N0_E2[1] <= N0_E1[0];    N2_E4[1] <= N2_E3[0];   N4_E6[1] <= N4_E5[0];   N6_S0[1] <= N6_E7[0];   E0_S2[1] <= E0_S1[0];   E3_S4[1] <= E3_S3[0];   E6_S6[1] <= E6_S5[0]; S4_W0[1] <= S3_W7[0];
	N0_E2[0] <= N0_E2[1];    N2_E4[0] <= N2_E4[1];   N4_E6[0] <= N4_E6[1];   N6_S0[0] <= N6_S0[1];   E0_S2[0] <= E0_S2[1];   E3_S4[0] <= E3_S4[1];   E6_S6[0] <= E6_S6[1]; S4_W0[0] <= S4_W0[1];
	N0_E3[1] <= N0_E2[0];    N2_E5[1] <= N2_E4[0];   N4_E7[1] <= N4_E6[0];   N6_S1[1] <= N6_S0[0];   E0_S3[1] <= E0_S2[0];   E3_S5[1] <= E3_S4[0];   E6_S7[1] <= E6_S6[0]; S4_W1[1] <= S4_W0[0];
	N0_E3[0] <= N0_E3[1];    N2_E5[0] <= N2_E5[1];   N4_E7[0] <= N4_E7[1];   N6_S1[0] <= N6_S1[1];   E0_S3[0] <= E0_S3[1];   E3_S5[0] <= E3_S5[1];   E6_S7[0] <= E6_S7[1]; S4_W1[0] <= S4_W1[1];
	N0_E4[1] <= N0_E3[0];    N2_E6[1] <= N2_E5[0];   N4_S0[1] <= N4_E7[0];   N6_S2[1] <= N6_S1[0];   E0_S4[1] <= E0_S3[0];   E3_S6[1] <= E3_S5[0];   E7_W0[1] <= E6_S7[0]; S4_W2[1] <= S4_W1[0];
	N0_E4[0] <= N0_E4[1];    N2_E6[0] <= N2_E6[1];   N4_S0[0] <= N4_S0[1];   N6_S2[0] <= N6_S2[1];   E0_S4[0] <= E0_S4[1];   E3_S6[0] <= E3_S6[1];   E7_W0[0] <= E7_W0[1]; S4_W2[0] <= S4_W2[1];
	N0_E5[1] <= N0_E4[0];    N2_E7[1] <= N2_E6[0];   N4_S1[1] <= N4_S0[0];   N6_S3[1] <= N6_S2[0];   E0_S5[1] <= E0_S4[0];   E3_S7[1] <= E3_S6[0];   E7_W1[1] <= E7_W0[0]; S4_W3[1] <= S4_W2[0];
	N0_E5[0] <= N0_E5[1];    N2_E7[0] <= N2_E7[1];   N4_S1[0] <= N4_S1[1];   N6_S3[0] <= N6_S3[1];   E0_S5[0] <= E0_S5[1];   E3_S7[0] <= E3_S7[1];   E7_W1[0] <= E7_W1[1]; S4_W3[0] <= S4_W3[1];
	N0_E6[1] <= N0_E5[0];    N2_S0[1] <= N2_E7[0];   N4_S2[1] <= N4_S1[0];   N6_S4[1] <= N6_S3[0];   E0_S6[1] <= E0_S5[0];   E4_W0[1] <= E3_S7[0];   E7_W2[1] <= E7_W1[0]; S4_W4[1] <= S4_W3[0];
	N0_E6[0] <= N0_E6[1];    N2_S0[0] <= N2_S0[1];   N4_S2[0] <= N4_S2[1];   N6_S4[0] <= N6_S4[1];   E0_S6[0] <= E0_S6[1];   E4_W0[0] <= E4_W0[1];   E7_W2[0] <= E7_W2[1]; S4_W4[0] <= S4_W4[1];
	N0_E7[1] <= N0_E6[0];    N2_S1[1] <= N2_S0[0];   N4_S3[1] <= N4_S2[0];   N6_S5[1] <= N6_S4[0];   E0_S7[1] <= E0_S6[0];   E4_W1[1] <= E4_W0[0];   E7_W3[1] <= E7_W2[0]; S4_W5[1] <= S4_W4[0];
	N0_E7[0] <= N0_E7[1];    N2_S1[0] <= N2_S1[1];   N4_S3[0] <= N4_S3[1];   N6_S5[0] <= N6_S5[1];   E0_S7[0] <= E0_S7[1];   E4_W1[0] <= E4_W1[1];   E7_W3[0] <= E7_W3[1]; S4_W5[0] <= S4_W5[1];
	N0_S0[1] <= N0_E7[0];    N2_S2[1] <= N2_S1[0];   N4_S4[1] <= N4_S3[0];   N6_S6[1] <= N6_S5[0];   E1_W0[1] <= E0_S7[0];   E4_W2[1] <= E4_W1[0];   E7_W4[1] <= E7_W3[0]; S4_W6[1] <= S4_W5[0];
	N0_S0[0] <= N0_S0[1];    N2_S2[0] <= N2_S2[1];   N4_S4[0] <= N4_S4[1];   N6_S6[0] <= N6_S6[1];   E1_W0[0] <= E1_W0[1];   E4_W2[0] <= E4_W2[1];   E7_W4[0] <= E7_W4[1]; S4_W6[0] <= S4_W6[1];
	N0_S1[1] <= N0_S0[0];    N2_S3[1] <= N2_S2[0];   N4_S5[1] <= N4_S4[0];   N6_S7[1] <= N6_S6[0];   E1_W1[1] <= E1_W0[0];   E4_W3[1] <= E4_W2[0];   E7_W5[1] <= E7_W4[0]; S4_W7[1] <= S4_W6[0];
	N0_S1[0] <= N0_S1[1];    N2_S3[0] <= N2_S3[1];   N4_S5[0] <= N4_S5[1];   N6_S7[0] <= N6_S7[1];   E1_W1[0] <= E1_W1[1];   E4_W3[0] <= E4_W3[1];   E7_W5[0] <= E7_W5[1]; S4_W7[0] <= S4_W7[1];
	N0_S2[1] <= N0_S1[0];    N2_S4[1] <= N2_S3[0];   N4_S6[1] <= N4_S5[0];   N6_W0[1] <= N6_S7[0];   E1_W2[1] <= E1_W1[0];   E4_W4[1] <= E4_W3[0];   E7_W6[1] <= E7_W5[0]; S5_W0[1] <= S4_W7[0];
	N0_S2[0] <= N0_S2[1];    N2_S4[0] <= N2_S4[1];   N4_S6[0] <= N4_S6[1];   N6_W0[0] <= N6_W0[1];   E1_W2[0] <= E1_W2[1];   E4_W4[0] <= E4_W4[1];   E7_W6[0] <= E7_W6[1]; S5_W0[0] <= S5_W0[1];
	N0_S3[1] <= N0_S2[0];    N2_S5[1] <= N2_S4[0];   N4_S7[1] <= N4_S6[0];   N6_W1[1] <= N6_W0[0];   E1_W3[1] <= E1_W2[0];   E4_W5[1] <= E4_W4[0];   E7_W7[1] <= E7_W6[0]; S5_W1[1] <= S5_W0[0];
	N0_S3[0] <= N0_S3[1];    N2_S5[0] <= N2_S5[1];   N4_S7[0] <= N4_S7[1];   N6_W1[0] <= N6_W1[1];   E1_W3[0] <= E1_W3[1];   E4_W5[0] <= E4_W5[1];   E7_W7[0] <= E7_W7[1]; S5_W1[0] <= S5_W1[1];
	N0_S4[1] <= N0_S3[0];    N2_S6[1] <= N2_S5[0];   N4_W0[1] <= N4_S7[0];   N6_W2[1] <= N6_W1[0];   E1_W4[1] <= E1_W3[0];   E4_W6[1] <= E4_W5[0];   E7_S0[1] <= E7_W7[0]; S5_W2[1] <= S5_W1[0];
	N0_S4[0] <= N0_S4[1];    N2_S6[0] <= N2_S6[1];   N4_W0[0] <= N4_W0[1];   N6_W2[0] <= N6_W2[1];   E1_W4[0] <= E1_W4[1];   E4_W6[0] <= E4_W6[1];   E7_S0[0] <= E7_S0[1]; S5_W2[0] <= S5_W2[1];
	N0_S5[1] <= N0_S4[0];    N2_S7[1] <= N2_S6[0];   N4_W1[1] <= N4_W0[0];   N6_W3[1] <= N6_W2[0];   E1_W5[1] <= E1_W4[0];   E4_W7[1] <= E4_W6[0];   E7_S1[1] <= E7_S0[0]; S5_W3[1] <= S5_W2[0];
	N0_S5[0] <= N0_S5[1];    N2_S7[0] <= N2_S7[1];   N4_W1[0] <= N4_W1[1];   N6_W3[0] <= N6_W3[1];   E1_W5[0] <= E1_W5[1];   E4_W7[0] <= E4_W7[1];   E7_S1[0] <= E7_S1[1]; S5_W3[0] <= S5_W3[1];
	N0_S6[1] <= N0_S5[0];    N2_W0[1] <= N2_S7[0];   N4_W2[1] <= N4_W1[0];   N6_W4[1] <= N6_W3[0];   E1_W6[1] <= E1_W5[0];   E4_S0[1] <= E4_W7[0];   E7_S2[1] <= E7_S1[0]; S5_W4[1] <= S5_W3[0];
	N0_S6[0] <= N0_S6[1];    N2_W0[0] <= N2_W0[1];   N4_W2[0] <= N4_W2[1];   N6_W4[0] <= N6_W4[1];   E1_W6[0] <= E1_W6[1];   E4_S0[0] <= E4_S0[1];   E7_S2[0] <= E7_S2[1]; S5_W4[0] <= S5_W4[1];
	N0_S7[1] <= N0_S6[0];    N2_W1[1] <= N2_W0[0];   N4_W3[1] <= N4_W2[0];   N6_W5[1] <= N6_W4[0];   E1_W7[1] <= E1_W6[0];   E4_S1[1] <= E4_S0[0];   E7_S3[1] <= E7_S2[0]; S5_W5[1] <= S5_W4[0];
	N0_S7[0] <= N0_S7[1];    N2_W1[0] <= N2_W1[1];   N4_W3[0] <= N4_W3[1];   N6_W5[0] <= N6_W5[1];   E1_W7[0] <= E1_W7[1];   E4_S1[0] <= E4_S1[1];   E7_S3[0] <= E7_S3[1]; S5_W5[0] <= S5_W5[1];
	N0_W0[1] <= N0_S7[0];    N2_W2[1] <= N2_W1[0];   N4_W4[1] <= N4_W3[0];   N6_W6[1] <= N6_W5[0];   E1_S0[1] <= E1_W7[0];   E4_S2[1] <= E4_S1[0];   E7_S4[1] <= E7_S3[0]; S5_W6[1] <= S5_W5[0];
	N0_W0[0] <= N0_W0[1];    N2_W2[0] <= N2_W2[1];   N4_W4[0] <= N4_W4[1];   N6_W6[0] <= N6_W6[1];   E1_S0[0] <= E1_S0[1];   E4_S2[0] <= E4_S2[1];   E7_S4[0] <= E7_S4[1]; S5_W6[0] <= S5_W6[1];
	N0_W1[1] <= N0_W0[0];    N2_W3[1] <= N2_W2[0];   N4_W5[1] <= N4_W4[0];   N6_W7[1] <= N6_W6[0];   E1_S1[1] <= E1_S0[0];   E4_S3[1] <= E4_S2[0];   E7_S5[1] <= E7_S4[0]; S5_W7[1] <= S5_W6[0];
	N0_W1[0] <= N0_W1[1];    N2_W3[0] <= N2_W3[1];   N4_W5[0] <= N4_W5[1];   N6_W7[0] <= N6_W7[1];   E1_S1[0] <= E1_S1[1];   E4_S3[0] <= E4_S3[1];   E7_S5[0] <= E7_S5[1]; S5_W7[0] <= S5_W7[1];
	N0_W2[1] <= N0_W1[0];    N2_W4[1] <= N2_W3[0];   N4_W6[1] <= N4_W5[0];   N7_E0[1] <= N6_W7[0];   E1_S2[1] <= E1_S1[0];   E4_S4[1] <= E4_S3[0];   E7_S6[1] <= E7_S5[0]; S6_W0[1] <= S5_W7[0];
	N0_W2[0] <= N0_W2[1];    N2_W4[0] <= N2_W4[1];   N4_W6[0] <= N4_W6[1];   N7_E0[0] <= N7_E0[1];   E1_S2[0] <= E1_S2[1];   E4_S4[0] <= E4_S4[1];   E7_S6[0] <= E7_S6[1]; S6_W0[0] <= S6_W0[1];
	N0_W3[1] <= N0_W2[0];    N2_W5[1] <= N2_W4[0];   N4_W7[1] <= N4_W6[0];   N7_E1[1] <= N7_E0[0];   E1_S3[1] <= E1_S2[0];   E4_S5[1] <= E4_S4[0];   E7_S7[1] <= E7_S6[0]; S6_W1[1] <= S6_W0[0];
	N0_W3[0] <= N0_W3[1];    N2_W5[0] <= N2_W5[1];   N4_W7[0] <= N4_W7[1];   N7_E1[0] <= N7_E1[1];   E1_S3[0] <= E1_S3[1];   E4_S5[0] <= E4_S5[1];   E7_S7[0] <= E7_S7[1]; S6_W1[0] <= S6_W1[1];
	N0_W4[1] <= N0_W3[0];    N2_W6[1] <= N2_W5[0];   N5_E0[1] <= N4_W7[0];   N7_E2[1] <= N7_E1[0];   E1_S4[1] <= E1_S3[0];   E4_S6[1] <= E4_S5[0];   S0_W0[1] <= E7_S7[0]; S6_W2[1] <= S6_W1[0];
	N0_W4[0] <= N0_W4[1];    N2_W6[0] <= N2_W6[1];   N5_E0[0] <= N5_E0[1];   N7_E2[0] <= N7_E2[1];   E1_S4[0] <= E1_S4[1];   E4_S6[0] <= E4_S6[1];   S0_W0[0] <= S0_W0[1]; S6_W2[0] <= S6_W2[1];
	N0_W5[1] <= N0_W4[0];    N2_W7[1] <= N2_W6[0];   N5_E1[1] <= N5_E0[0];   N7_E3[1] <= N7_E2[0];   E1_S5[1] <= E1_S4[0];   E4_S7[1] <= E4_S6[0];   S0_W1[1] <= S0_W0[0]; S6_W3[1] <= S6_W2[0];
	N0_W5[0] <= N0_W5[1];    N2_W7[0] <= N2_W7[1];   N5_E1[0] <= N5_E1[1];   N7_E3[0] <= N7_E3[1];   E1_S5[0] <= E1_S5[1];   E4_S7[0] <= E4_S7[1];   S0_W1[0] <= S0_W1[1]; S6_W3[0] <= S6_W3[1];
	N0_W6[1] <= N0_W5[0];    N3_E0[1] <= N2_W7[0];   N5_E2[1] <= N5_E1[0];   N7_E4[1] <= N7_E3[0];   E1_S6[1] <= E1_S5[0];   E5_W0[1] <= E4_S7[0];   S0_W2[1] <= S0_W1[0]; S6_W4[1] <= S6_W3[0];
	N0_W6[0] <= N0_W6[1];    N3_E0[0] <= N3_E0[1];   N5_E2[0] <= N5_E2[1];   N7_E4[0] <= N7_E4[1];   E1_S6[0] <= E1_S6[1];   E5_W0[0] <= E5_W0[1];   S0_W2[0] <= S0_W2[1]; S6_W4[0] <= S6_W4[1];
	N0_W7[1] <= N0_W6[0];    N3_E1[1] <= N3_E0[0];   N5_E3[1] <= N5_E2[0];   N7_E5[1] <= N7_E4[0];   E1_S7[1] <= E1_S6[0];   E5_W1[1] <= E5_W0[0];   S0_W3[1] <= S0_W2[0]; S6_W5[1] <= S6_W4[0];
	N0_W7[0] <= N0_W7[1];    N3_E1[0] <= N3_E1[1];   N5_E3[0] <= N5_E3[1];   N7_E5[0] <= N7_E5[1];   E1_S7[0] <= E1_S7[1];   E5_W1[0] <= E5_W1[1];   S0_W3[0] <= S0_W3[1]; S6_W5[0] <= S6_W5[1];
	N1_E0[1] <= N0_W7[0];    N3_E2[1] <= N3_E1[0];   N5_E4[1] <= N5_E3[0];   N7_E6[1] <= N7_E5[0];   E2_W0[1] <= E1_S7[0];   E5_W2[1] <= E5_W1[0];   S0_W4[1] <= S0_W3[0]; S6_W6[1] <= S6_W5[0];
	N1_E0[0] <= N1_E0[1];    N3_E2[0] <= N3_E2[1];   N5_E4[0] <= N5_E4[1];   N7_E6[0] <= N7_E6[1];   E2_W0[0] <= E2_W0[1];   E5_W2[0] <= E5_W2[1];   S0_W4[0] <= S0_W4[1]; S6_W6[0] <= S6_W6[1];
	N1_E1[1] <= N1_E0[0];    N3_E3[1] <= N3_E2[0];   N5_E5[1] <= N5_E4[0];   N7_E7[1] <= N7_E6[0];   E2_W1[1] <= E2_W0[0];   E5_W3[1] <= E5_W2[0];   S0_W5[1] <= S0_W4[0]; S6_W7[1] <= S6_W6[0];
	N1_E1[0] <= N1_E1[1];    N3_E3[0] <= N3_E3[1];   N5_E5[0] <= N5_E5[1];   N7_E7[0] <= N7_E7[1];   E2_W1[0] <= E2_W1[1];   E5_W3[0] <= E5_W3[1];   S0_W5[0] <= S0_W5[1]; S6_W7[0] <= S6_W7[1];
	N1_E2[1] <= N1_E1[0];    N3_E4[1] <= N3_E3[0];   N5_E6[1] <= N5_E5[0];   N7_S0[1] <= N7_E7[0];   E2_W2[1] <= E2_W1[0];   E5_W4[1] <= E5_W3[0];   S0_W6[1] <= S0_W5[0]; S7_W0[1] <= S6_W7[0];
	N1_E2[0] <= N1_E2[1];    N3_E4[0] <= N3_E4[1];   N5_E6[0] <= N5_E6[1];   N7_S0[0] <= N7_S0[1];   E2_W2[0] <= E2_W2[1];   E5_W4[0] <= E5_W4[1];   S0_W6[0] <= S0_W6[1]; S7_W0[0] <= S7_W0[1];
	N1_E3[1] <= N1_E2[0];    N3_E5[1] <= N3_E4[0];   N5_E7[1] <= N5_E6[0];   N7_S1[1] <= N7_S0[0];   E2_W3[1] <= E2_W2[0];   E5_W5[1] <= E5_W4[0];   S0_W7[1] <= S0_W6[0]; S7_W1[1] <= S7_W0[0];
	N1_E3[0] <= N1_E3[1];    N3_E5[0] <= N3_E5[1];   N5_E7[0] <= N5_E7[1];   N7_S1[0] <= N7_S1[1];   E2_W3[0] <= E2_W3[1];   E5_W5[0] <= E5_W5[1];   S0_W7[0] <= S0_W7[1]; S7_W1[0] <= S7_W1[1];
	N1_E4[1] <= N1_E3[0];    N3_E6[1] <= N3_E5[0];   N5_S0[1] <= N5_E7[0];   N7_S2[1] <= N7_S1[0];   E2_W4[1] <= E2_W3[0];   E5_W6[1] <= E5_W5[0];   S1_W0[1] <= S0_W7[0]; S7_W2[1] <= S7_W1[0];
	N1_E4[0] <= N1_E4[1];    N3_E6[0] <= N3_E6[1];   N5_S0[0] <= N5_S0[1];   N7_S2[0] <= N7_S2[1];   E2_W4[0] <= E2_W4[1];   E5_W6[0] <= E5_W6[1];   S1_W0[0] <= S1_W0[1]; S7_W2[0] <= S7_W2[1];
	N1_E5[1] <= N1_E4[0];    N3_E7[1] <= N3_E6[0];   N5_S1[1] <= N5_S0[0];   N7_S3[1] <= N7_S2[0];   E2_W5[1] <= E2_W4[0];   E5_W7[1] <= E5_W6[0];   S1_W1[1] <= S1_W0[0]; S7_W3[1] <= S7_W2[0];
	N1_E5[0] <= N1_E5[1];    N3_E7[0] <= N3_E7[1];   N5_S1[0] <= N5_S1[1];   N7_S3[0] <= N7_S3[1];   E2_W5[0] <= E2_W5[1];   E5_W7[0] <= E5_W7[1];   S1_W1[0] <= S1_W1[1]; S7_W3[0] <= S7_W3[1];
	N1_E6[1] <= N1_E5[0];    N3_S0[1] <= N3_E7[0];   N5_S2[1] <= N5_S1[0];   N7_S4[1] <= N7_S3[0];   E2_W6[1] <= E2_W5[0];   E5_S0[1] <= E5_W7[0];   S1_W2[1] <= S1_W1[0]; S7_W4[1] <= S7_W3[0];
	N1_E6[0] <= N1_E6[1];    N3_S0[0] <= N3_S0[1];   N5_S2[0] <= N5_S2[1];   N7_S4[0] <= N7_S4[1];   E2_W6[0] <= E2_W6[1];   E5_S0[0] <= E5_S0[1];   S1_W2[0] <= S1_W2[1]; S7_W4[0] <= S7_W4[1];
	N1_E7[1] <= N1_E6[0];    N3_S1[1] <= N3_S0[0];   N5_S3[1] <= N5_S2[0];   N7_S5[1] <= N7_S4[0];   E2_W7[1] <= E2_W6[0];   E5_S1[1] <= E5_S0[0];   S1_W3[1] <= S1_W2[0]; S7_W5[1] <= S7_W4[0];
	N1_E7[0] <= N1_E7[1];    N3_S1[0] <= N3_S1[1];   N5_S3[0] <= N5_S3[1];   N7_S5[0] <= N7_S5[1];   E2_W7[0] <= E2_W7[1];   E5_S1[0] <= E5_S1[1];   S1_W3[0] <= S1_W3[1]; S7_W5[0] <= S7_W5[1];
	N1_S0[1] <= N1_E7[0];    N3_S2[1] <= N3_S1[0];   N5_S4[1] <= N5_S3[0];   N7_S6[1] <= N7_S5[0];   E2_S0[1] <= E2_W7[0];   E5_S2[1] <= E5_S1[0];   S1_W4[1] <= S1_W3[0]; S7_W6[1] <= S7_W5[0];
	N1_S0[0] <= N1_S0[1];    N3_S2[0] <= N3_S2[1];   N5_S4[0] <= N5_S4[1];   N7_S6[0] <= N7_S6[1];   E2_S0[0] <= E2_S0[1];   E5_S2[0] <= E5_S2[1];   S1_W4[0] <= S1_W4[1]; S7_W6[0] <= S7_W6[1];
	N1_S1[1] <= N1_S0[0];    N3_S3[1] <= N3_S2[0];   N5_S5[1] <= N5_S4[0];   N7_S7[1] <= N7_S6[0];   E2_S1[1] <= E2_S0[0];   E5_S3[1] <= E5_S2[0];   S1_W5[1] <= S1_W4[0]; S7_W7[1] <= S7_W6[0];
	N1_S1[0] <= N1_S1[1];    N3_S3[0] <= N3_S3[1];   N5_S5[0] <= N5_S5[1];   N7_S7[0] <= N7_S7[1];   E2_S1[0] <= E2_S1[1];   E5_S3[0] <= E5_S3[1];   S1_W5[0] <= S1_W5[1]; S7_W7[0] <= S7_W7[1];
	N1_S2[1] <= N1_S1[0];    N3_S4[1] <= N3_S3[0];   N5_S6[1] <= N5_S5[0];   N7_W0[1] <= N7_S7[0];   E2_S2[1] <= E2_S1[0];   E5_S4[1] <= E5_S3[0];   S1_W6[1] <= S1_W5[0];                  
	N1_S2[0] <= N1_S2[1];    N3_S4[0] <= N3_S4[1];   N5_S6[0] <= N5_S6[1];   N7_W0[0] <= N7_W0[1];   E2_S2[0] <= E2_S2[1];   E5_S4[0] <= E5_S4[1];   S1_W6[0] <= S1_W6[1];                  
	N1_S3[1] <= N1_S2[0];    N3_S5[1] <= N3_S4[0];   N5_S7[1] <= N5_S6[0];   N7_W1[1] <= N7_W0[0];   E2_S3[1] <= E2_S2[0];   E5_S5[1] <= E5_S4[0];   S1_W7[1] <= S1_W6[0];                  
	N1_S3[0] <= N1_S3[1];    N3_S5[0] <= N3_S5[1];   N5_S7[0] <= N5_S7[1];   N7_W1[0] <= N7_W1[1];   E2_S3[0] <= E2_S3[1];   E5_S5[0] <= E5_S5[1];   S1_W7[0] <= S1_W7[1];                  
	N1_S4[1] <= N1_S3[0];    N3_S6[1] <= N3_S5[0];   N5_W0[1] <= N5_S7[0];   N7_W2[1] <= N7_W1[0];   E2_S4[1] <= E2_S3[0];   E5_S6[1] <= E5_S5[0];   S2_W0[1] <= S1_W7[0];                  
	N1_S4[0] <= N1_S4[1];    N3_S6[0] <= N3_S6[1];   N5_W0[0] <= N5_W0[1];   N7_W2[0] <= N7_W2[1];   E2_S4[0] <= E2_S4[1];   E5_S6[0] <= E5_S6[1];   S2_W0[0] <= S2_W0[1];                  
	N1_S5[1] <= N1_S4[0];    N3_S7[1] <= N3_S6[0];   N5_W1[1] <= N5_W0[0];   N7_W3[1] <= N7_W2[0];   E2_S5[1] <= E2_S4[0];   E5_S7[1] <= E5_S6[0];   S2_W1[1] <= S2_W0[0];                  
	N1_S5[0] <= N1_S5[1];    N3_S7[0] <= N3_S7[1];   N5_W1[0] <= N5_W1[1];   N7_W3[0] <= N7_W3[1];   E2_S5[0] <= E2_S5[1];   E5_S7[0] <= E5_S7[1];   S2_W1[0] <= S2_W1[1];                  
	N1_S6[1] <= N1_S5[0];    N3_W0[1] <= N3_S7[0];   N5_W2[1] <= N5_W1[0];   N7_W4[1] <= N7_W3[0];   E2_S6[1] <= E2_S5[0];   E6_W0[1] <= E5_S7[0];   S2_W2[1] <= S2_W1[0];                  
	N1_S6[0] <= N1_S6[1];    N3_W0[0] <= N3_W0[1];   N5_W2[0] <= N5_W2[1];   N7_W4[0] <= N7_W4[1];   E2_S6[0] <= E2_S6[1];   E6_W0[0] <= E6_W0[1];   S2_W2[0] <= S2_W2[1];                  
	N1_S7[1] <= N1_S6[0];    N3_W1[1] <= N3_W0[0];   N5_W3[1] <= N5_W2[0];   N7_W5[1] <= N7_W4[0];   E2_S7[1] <= E2_S6[0];   E6_W1[1] <= E6_W0[0];   S2_W3[1] <= S2_W2[0];                  
	N1_S7[0] <= N1_S7[1];    N3_W1[0] <= N3_W1[1];   N5_W3[0] <= N5_W3[1];   N7_W5[0] <= N7_W5[1];   E2_S7[0] <= E2_S7[1];   E6_W1[0] <= E6_W1[1];   S2_W3[0] <= S2_W3[1];                  
	N1_W0[1] <= N1_S7[0];    N3_W2[1] <= N3_W1[0];   N5_W4[1] <= N5_W3[0];   N7_W6[1] <= N7_W5[0];   E3_W0[1] <= E2_S7[0];   E6_W2[1] <= E6_W1[0];   S2_W4[1] <= S2_W3[0];                  
	N1_W0[0] <= N1_W0[1];    N3_W2[0] <= N3_W2[1];   N5_W4[0] <= N5_W4[1];   N7_W6[0] <= N7_W6[1];   E3_W0[0] <= E3_W0[1];   E6_W2[0] <= E6_W2[1];   S2_W4[0] <= S2_W4[1];                  
	N1_W1[1] <= N1_W0[0];    N3_W3[1] <= N3_W2[0];   N5_W5[1] <= N5_W4[0];   N7_W7[1] <= N7_W6[0];   E3_W1[1] <= E3_W0[0];   E6_W3[1] <= E6_W2[0];   S2_W5[1] <= S2_W4[0];                  
	N1_W1[0] <= N1_W1[1];    N3_W3[0] <= N3_W3[1];   N5_W5[0] <= N5_W5[1];   N7_W7[0] <= N7_W7[1];   E3_W1[0] <= E3_W1[1];   E6_W3[0] <= E6_W3[1];   S2_W5[0] <= S2_W5[1];                  
	N1_W2[1] <= N1_W1[0];    N3_W4[1] <= N3_W3[0];   N5_W6[1] <= N5_W5[0];   E0_W0[1] <= N7_W7[0];   E3_W2[1] <= E3_W1[0];   E6_W4[1] <= E6_W3[0];   S2_W6[1] <= S2_W5[0];                  
	N1_W2[0] <= N1_W2[1];    N3_W4[0] <= N3_W4[1];   N5_W6[0] <= N5_W6[1];   E0_W0[0] <= E0_W0[1];   E3_W2[0] <= E3_W2[1];   E6_W4[0] <= E6_W4[1];   S2_W6[0] <= S2_W6[1];                  
	N1_W3[1] <= N1_W2[0];    N3_W5[1] <= N3_W4[0];   N5_W7[1] <= N5_W6[0];   E0_W1[1] <= E0_W0[0];   E3_W3[1] <= E3_W2[0];   E6_W5[1] <= E6_W4[0];   S2_W7[1] <= S2_W6[0];                  
	N1_W3[0] <= N1_W3[1];    N3_W5[0] <= N3_W5[1];   N5_W7[0] <= N5_W7[1];   E0_W1[0] <= E0_W1[1];   E3_W3[0] <= E3_W3[1];   E6_W5[0] <= E6_W5[1];   S2_W7[0] <= S2_W7[1];                  
	N1_W4[1] <= N1_W3[0];    N3_W6[1] <= N3_W5[0];   N6_E0[1] <= N5_W7[0];   E0_W2[1] <= E0_W1[0];   E3_W4[1] <= E3_W3[0];   E6_W6[1] <= E6_W5[0];   S3_W0[1] <= S2_W7[0];                  
	N1_W4[0] <= N1_W4[1];    N3_W6[0] <= N3_W6[1];   N6_E0[0] <= N6_E0[1];   E0_W2[0] <= E0_W2[1];   E3_W4[0] <= E3_W4[1];   E6_W6[0] <= E6_W6[1];   S3_W0[0] <= S3_W0[1];                  
	N1_W5[1] <= N1_W4[0];    N3_W7[1] <= N3_W6[0];   N6_E1[1] <= N6_E0[0];   E0_W3[1] <= E0_W2[0];   E3_W5[1] <= E3_W4[0];   E6_W7[1] <= E6_W6[0];   S3_W1[1] <= S3_W0[0];                  
	N1_W5[0] <= N1_W5[1];    N3_W7[0] <= N3_W7[1];   N6_E1[0] <= N6_E1[1];   E0_W3[0] <= E0_W3[1];   E3_W5[0] <= E3_W5[1];   E6_W7[0] <= E6_W7[1];   S3_W1[0] <= S3_W1[1];                  
	N1_W6[1] <= N1_W5[0];    N4_E0[1] <= N3_W7[0];   N6_E2[1] <= N6_E1[0];   E0_W4[1] <= E0_W3[0];   E3_W6[1] <= E3_W5[0];   E6_S0[1] <= E6_W7[0];   S3_W2[1] <= S3_W1[0];                  
	N1_W6[0] <= N1_W6[1];    N4_E0[0] <= N4_E0[1];   N6_E2[0] <= N6_E2[1];   E0_W4[0] <= E0_W4[1];   E3_W6[0] <= E3_W6[1];   E6_S0[0] <= E6_S0[1];   S3_W2[0] <= S3_W2[1];                  
	N1_W7[1] <= N1_W6[0];    N4_E1[1] <= N4_E0[0];   N6_E3[1] <= N6_E2[0];   E0_W5[1] <= E0_W4[0];   E3_W7[1] <= E3_W6[0];   E6_S1[1] <= E6_S0[0];   S3_W3[1] <= S3_W2[0];                  
	N1_W7[0] <= N1_W7[1];    N4_E1[0] <= N4_E1[1];   N6_E3[0] <= N6_E3[1];   E0_W5[0] <= E0_W5[1];   E3_W7[0] <= E3_W7[1];   E6_S1[0] <= E6_S1[1];   S3_W3[0] <= S3_W3[1];                  
	N2_E0[1] <= N1_W7[0];    N4_E2[1] <= N4_E1[0];   N6_E4[1] <= N6_E3[0];   E0_W6[1] <= E0_W5[0];   E3_S0[1] <= E3_W7[0];   E6_S2[1] <= E6_S1[0];   S3_W4[1] <= S3_W3[0];                  
	N2_E0[0] <= N2_E0[1];    N4_E2[0] <= N4_E2[1];   N6_E4[0] <= N6_E4[1];   E0_W6[0] <= E0_W6[1];   E3_S0[0] <= E3_S0[1];   E6_S2[0] <= E6_S2[1];   S3_W4[0] <= S3_W4[1];                  
	N2_E1[1] <= N2_E0[0];    N4_E3[1] <= N4_E2[0];   N6_E5[1] <= N6_E4[0];   E0_W7[1] <= E0_W6[0];   E3_S1[1] <= E3_S0[0];   E6_S3[1] <= E6_S2[0];   S3_W5[1] <= S3_W4[0];                  
	N2_E1[0] <= N2_E1[1];    N4_E3[0] <= N4_E3[1];   N6_E5[0] <= N6_E5[1];   E0_W7[0] <= E0_W7[1];   E3_S1[0] <= E3_S1[1];   E6_S3[0] <= E6_S3[1];   S3_W5[0] <= S3_W5[1]; 
                 
                      
	

	end
	end
	end
	
	endmodule
		
