module FPGA_testbench();


reg [5119:0] CB_config_stream ;
reg [7423:0] CLB_config_stream;
reg [319:0] IO_config_stream;
reg [19199:0] SB_config_stream;

reg [7679:0] SB_config_stream0;
reg [7679:0] SB_config_stream1;
reg [3839:0] SB_config_stream2;


reg [5119:0] CB_config_stream_final ;
reg [7423:0] CLB_config_stream_final;
reg [319:0] IO_config_stream_final;
reg [19199:0] SB_config_stream_final;


wire cb_prgm_b_out,sb_prgm_b_out,io_prgm_b_out,CLB_prgm_b_out;
reg GWE;


wire G0,G1,G2,G3,G4,G5,G6,G7;
integer i0,i1,i2,k,l,m;


inout V00_0,V00_1,V00_2,V00_3,V00_4,V00_5,V00_6,V00_7,V01_0,V01_1,V01_2,V01_3,V01_4,V01_5,V01_6,V01_7,V02_0,V02_1,V02_2,V02_3,V02_4,V02_5,V02_6,V02_7,V03_0,V03_1,V03_2,V03_3,V03_4,V03_5,V03_6,V03_7,V04_0,V04_1,V04_2,V04_3,V04_4,V04_5,V04_6,V04_7,   
H10_0,H10_1,H10_2,H10_3,H10_4,H10_5,H10_6,H10_7,H11_0,H11_1,H11_2,H11_3,H11_4,H11_5,H11_6,H11_7,H20_0,H20_1,H20_2,H20_3,H20_4,H20_5,H20_6,H20_7,H21_0,H21_1,H21_2,H21_3,H21_4,H21_5,H21_6,H21_7,
H30_0,H30_1,H30_2,H30_3,H30_4,H30_5,H30_6,H30_7,H31_0,H31_1,H31_2,H31_3,H31_4,H31_5,H31_6,H31_7,H40_0,H40_1,H40_2,H40_3,H40_4,H40_5,H40_6,H40_7,H41_0,H41_1,H41_2,H41_3,H41_4,H41_5,H41_6,H41_7,
H50_3,H50_4,H50_5,H50_6,H50_7,H51_0,H51_1,H51_2,H51_3,H51_4,H51_5,H51_6,H51_7,
V60_0,V60_1,V60_2,V60_3,V60_4,V60_5,V60_6,V60_7,V61_0,V61_1,V61_2,V61_3,V61_4,V61_5,V61_6,V61_7,V62_0,V62_1,V62_2,V62_3,V62_4,V62_5,V62_6,V62_7,V63_0,V63_1,V63_2,V63_3,V63_4,V63_5,V63_6,V63_7,V64_0,V64_1,V64_2,V64_3,V64_4,V64_5,V64_6,V64_7;

reg V000,V001,V002,V003,V004,V005,V006,V007,V010,V011,V012,V013,V014,V015,V016,V017,V020,V021,V022,V023,V024,V025,V026,V027,V030,V031,V032,V033,V034,V035,V036,V037,V040,V041,V042,V043,V044,V045,V046,V047,   
H100,H101,H102,H103,H104,H105,H106,H107,H110,H111,H112,H113,H114,H115,H116,H117,H200,H201,H202,H203,H204,H205,H206,H207,H210,H211,H212,H213,H214,H215,H216,H217,
H300,H301,H302,H303,H304,H305,H306,H307,H310,H311,H312,H313,H314,H315,H316,H317,H400,H401,H402,H403,H404,H405,H406,H407,H410,H411,H412,H413,H414,H415,H416,H417,
H503,H504,H505,H506,H507,H510,H511,H512,H513,H514,H515,H516,H517,
V600,V601,V602,V603,V604,V605,V606,V607,V610,V611,V612,V613,V614,V615,V616,V617,V620,V621,V622,V623,V624,V625,V626,V627,V630,V631,V632,V633,V634,V635,V636,V637,V640,V641,V642,V643,V644,V645,V646,V647;

 
value v000(.in(V000) , .out(V00_0) );           value v600(.in(V600) , .out(V60_0) );
value v001(.in(V001) , .out(V00_1) );           value v601(.in(V601) , .out(V60_1) );
value v002(.in(V002) , .out(V00_2) );           value v602(.in(V602) , .out(V60_2) );
value v003(.in(V003) , .out(V00_3) );           value v603(.in(V603) , .out(V60_3) );
value v004(.in(V004) , .out(V00_4) );           value v604(.in(V604) , .out(V60_4) );
value v005(.in(V005) , .out(V00_5) );           value v605(.in(V605) , .out(V60_5) );
value v006(.in(V006) , .out(V00_6) );           value v606(.in(V606) , .out(V60_6) );
value v007(.in(V007) , .out(V00_7) );           value v607(.in(V607) , .out(V60_7) );
                                                
value v010(.in(V010) , .out(V01_0) );           value v610(.in(V610) , .out(V61_0) );
value v011(.in(V011) , .out(V01_1) );           value v611(.in(V611) , .out(V61_1) );
value v012(.in(V012) , .out(V01_2) );           value v612(.in(V612) , .out(V61_2) );
value v013(.in(V013) , .out(V01_3) );           value v613(.in(V613) , .out(V61_3) );
value v014(.in(V014) , .out(V01_4) );           value v614(.in(V614) , .out(V61_4) );
value v015(.in(V015) , .out(V01_5) );           value v615(.in(V615) , .out(V61_5) );
value v016(.in(V016) , .out(V01_6) );           value v616(.in(V616) , .out(V61_6) );
value v017(.in(V017) , .out(V01_7) );           value v617(.in(V617) , .out(V61_7) );
                                                
value v020(.in(V020) , .out(V02_0) );           value v620(.in(V620) , .out(V62_0) );
value v021(.in(V021) , .out(V02_1) );           value v621(.in(V621) , .out(V62_1) );
value v022(.in(V022) , .out(V02_2) );           value v622(.in(V622) , .out(V62_2) );
value v023(.in(V023) , .out(V02_3) );           value v623(.in(V623) , .out(V62_3) );
value v024(.in(V024) , .out(V02_4) );           value v624(.in(V624) , .out(V62_4) );
value v025(.in(V025) , .out(V02_5) );           value v625(.in(V625) , .out(V62_5) );
value v026(.in(V026) , .out(V02_6) );           value v626(.in(V626) , .out(V62_6) );
value v027(.in(V027) , .out(V02_7) );           value v627(.in(V627) , .out(V62_7) );
                                                
value v030(.in(V030) , .out(V03_0) );           value v630(.in(V630) , .out(V63_0) );
value v031(.in(V031) , .out(V03_1) );           value v631(.in(V631) , .out(V63_1) );
value v032(.in(V032) , .out(V03_2) );           value v632(.in(V632) , .out(V63_2) );
value v033(.in(V033) , .out(V03_3) );           value v633(.in(V633) , .out(V63_3) );
value v034(.in(V034) , .out(V03_4) );           value v634(.in(V634) , .out(V63_4) );
value v035(.in(V035) , .out(V03_5) );           value v635(.in(V635) , .out(V63_5) );
value v036(.in(V036) , .out(V03_6) );           value v636(.in(V636) , .out(V63_6) );
value v037(.in(V037) , .out(V03_7) );           value v637(.in(V637) , .out(V63_7) );
                                                
value v040(.in(V040) , .out(V04_0) );           value v640(.in(V640) , .out(V64_0) );
value v041(.in(V041) , .out(V04_1) );           value v641(.in(V641) , .out(V64_1) );
value v042(.in(V042) , .out(V04_2) );           value v642(.in(V642) , .out(V64_2) );
value v043(.in(V043) , .out(V04_3) );           value v643(.in(V643) , .out(V64_3) );
value v044(.in(V044) , .out(V04_4) );           value v644(.in(V644) , .out(V64_4) );
value v045(.in(V045) , .out(V04_5) );           value v645(.in(V645) , .out(V64_5) );
value v046(.in(V046) , .out(V04_6) );           value v646(.in(V646) , .out(V64_6) );
value v047(.in(V047) , .out(V04_7) );           value v647(.in(V647) , .out(V64_7) );

value h100(.in(H100) , .out(H10_0) );           value h200(.in(H200) , .out(H20_0) );
value h101(.in(H101) , .out(H10_1) );           value h201(.in(H201) , .out(H20_1) );
value h102(.in(H102) , .out(H10_2) );           value h202(.in(H202) , .out(H20_2) );
value h103(.in(H103) , .out(H10_3) );           value h203(.in(H203) , .out(H20_3) );
value h104(.in(H104) , .out(H10_4) );           value h204(.in(H204) , .out(H20_4) );
value h105(.in(H105) , .out(H10_5) );           value h205(.in(H205) , .out(H20_5) );
value h106(.in(H106) , .out(H10_6) );           value h206(.in(H206) , .out(H20_6) );
value h107(.in(H107) , .out(H10_7) );           value h207(.in(H207) , .out(H20_7) );
                                                
value h110(.in(H110) , .out(H11_0) );           value h210(.in(H210) , .out(H21_0) );
value h111(.in(H111) , .out(H11_1) );           value h211(.in(H211) , .out(H21_1) );
value h112(.in(H112) , .out(H11_2) );           value h212(.in(H212) , .out(H21_2) );
value h113(.in(H113) , .out(H11_3) );           value h213(.in(H213) , .out(H21_3) );
value h114(.in(H114) , .out(H11_4) );           value h214(.in(H214) , .out(H21_4) );
value h115(.in(H115) , .out(H11_5) );           value h215(.in(H215) , .out(H21_5) );
value h116(.in(H116) , .out(H11_6) );           value h216(.in(H216) , .out(H21_6) );
value h117(.in(H117) , .out(H11_7) );           value h217(.in(H217) , .out(H21_7) );

value h300(.in(H300) , .out(H30_0) );           value h400(.in(H400) , .out(H40_0) );
value h301(.in(H301) , .out(H30_1) );           value h401(.in(H401) , .out(H40_1) );
value h302(.in(H302) , .out(H30_2) );           value h402(.in(H402) , .out(H40_2) );
value h303(.in(H303) , .out(H30_3) );           value h403(.in(H403) , .out(H40_3) );
value h304(.in(H304) , .out(H30_4) );           value h404(.in(H404) , .out(H40_4) );
value h305(.in(H305) , .out(H30_5) );           value h405(.in(H405) , .out(H40_5) );
value h306(.in(H306) , .out(H30_6) );           value h406(.in(H406) , .out(H40_6) );
value h307(.in(H307) , .out(H30_7) );           value h407(.in(H407) , .out(H40_7) );
                                                
value h310(.in(H310) , .out(H31_0) );           value h410(.in(H410) , .out(H41_0) );
value h311(.in(H311) , .out(H31_1) );           value h411(.in(H411) , .out(H41_1) );
value h312(.in(H312) , .out(H31_2) );           value h412(.in(H412) , .out(H41_2) );
value h313(.in(H313) , .out(H31_3) );           value h413(.in(H413) , .out(H41_3) );
value h314(.in(H314) , .out(H31_4) );           value h414(.in(H414) , .out(H41_4) );
value h315(.in(H315) , .out(H31_5) );           value h415(.in(H415) , .out(H41_5) );
value h316(.in(H316) , .out(H31_6) );           value h416(.in(H416) , .out(H41_6) );
value h317(.in(H317) , .out(H31_7) );           value h417(.in(H417) , .out(H41_7) );

value h500(.in(H500) , .out(H50_0) );           value h510(.in(H510) , .out(H51_0) );
value h501(.in(H501) , .out(H50_1) );           value h511(.in(H511) , .out(H51_1) );
value h502(.in(H502) , .out(H50_2) );           value h512(.in(H512) , .out(H51_2) );
value h503(.in(H503) , .out(H50_3) );           value h513(.in(H513) , .out(H51_3) );
value h504(.in(H504) , .out(H50_4) );           value h514(.in(H514) , .out(H51_4) );
value h505(.in(H505) , .out(H50_5) );           value h515(.in(H515) , .out(H51_5) );
value h506(.in(H506) , .out(H50_6) );           value h516(.in(H516) , .out(H51_6) );
value h507(.in(H507) , .out(H50_7) );           value h517(.in(H517) , .out(H51_7) );      

reg clk,reset,prgm_b,CLB_prgm_b,cb_prgm_b,sb_prgm_b,bit_in_CLB,bit_in_CB,bit_in_SB,bit_in_SB_2,sb_prgm_b_in,
cb_prgm_b_in,CLB_prgm_b_in,sb_prgm_b_2,io_prgm_b_in,bit_in_IO,io_prgm_b;

integer CB_count,SB_count,IO_count,CLB_count,CLB_counter,CB_counter,SB_counter,IO_counter;


FPGA FPGA4x4(.V00_0(V00_0),.V00_1(V00_1),.V00_2(V00_2),.V00_3(V00_3),.V00_4(V00_4),.V00_5(V00_5),.V00_6(V00_6),.V00_7(V00_7),.V01_0(V01_0),
.V01_1(V01_1),.V01_2(V01_2),.V01_3(V01_3),.V01_4(V01_4),.V01_5(V01_5),.V01_6(V01_6),.V01_7(V01_7),.V02_0(V02_0),.V02_1(V02_1),.V02_2(V02_2),
.V02_3(V02_3),.V02_4(V02_4),.V02_5(V02_5),.V02_6(V02_6),.V02_7(V02_7),.V03_0(V03_0),.V03_1(V03_1),.V03_2(V03_2),.V03_3(V03_3),.V03_4(V03_4),
.V03_5(V03_5),.V03_6(V03_6),.V03_7(V03_7),.V04_0(V04_0),.V04_1(V04_1),.V04_2(V04_2),.V04_3(V04_3),.V04_4(V04_4),.V04_5(V04_5),.V04_6(V04_6),.V04_7(V04_7),.H10_0(H10_0),.H10_1(H10_1),.H10_2(H10_2),.H10_3(H10_3),.H10_4(H10_4),.H10_5(H10_5),.H10_6(H10_6),.H10_7(H10_7),.H11_0(H11_0),.H11_1(H11_1),
.H11_2(H11_2),.H11_3(H11_3),.H11_4(H11_4),.H11_5(H11_5),.H11_6(H11_6),.H11_7(H11_7),
.H20_0(H20_0),.H20_1(H20_1),.H20_2(H20_2),.H20_3(H20_3),.H20_4(H20_4),.H20_5(H20_5),.H20_6(H20_6),.H20_7(H20_7),.H21_0(H21_0),.H21_1(H21_1),
.H21_2(H21_2),.H21_3(H21_3),.H21_4(H21_4),.H21_5(H21_5),.H21_6(H21_6),.H21_7(H21_7),
      .H30_0(H30_0),.H30_1(H30_1),.H30_2(H30_2),.H30_3(H30_3),.H30_4(H30_4),.H30_5(H30_5),.H30_6(H30_6),.H30_7(H30_7),.H31_0(H31_0),.H31_1(H31_1),
.H31_2(H31_2),.H31_3(H31_3),.H31_4(H31_4),.H31_5(H31_5),.H31_6(H31_6),.H31_7(H31_7),
      .H40_0(H40_0),.H40_1(H40_1),.H40_2(H40_2),.H40_3(H40_3),.H40_4(H40_4),.H40_5(H40_5),.H40_6(H40_6),.H40_7(H40_7),.H41_0(H41_0),.H41_1(H41_1),
.H41_2(H41_2),.H41_3(H41_3),.H41_4(H41_4),.H41_5(H41_5),.H41_6(H41_6),.H41_7(H41_7),
	  .H50_0(H50_0),.H50_1(H50_1),.H50_2(H50_2),.H50_3(H50_3),.H50_4(H50_4),.H50_5(H50_5),.H50_6(H50_6),.H50_7(H50_7),.H51_0(H51_0),.H51_1(H51_1),
.H51_2(H51_2),.H51_3(H51_3),.H51_4(H51_4),.H51_5(H51_5),.H51_6(H51_6),.H51_7(H51_7),
       .V60_0(V60_0),.V60_1(V60_1),.V60_2(V60_2),.V60_3(V60_3),.V60_4(V60_4),.V60_5(V60_5),.V60_6(V60_6),.V60_7(V60_7),.V61_0(V61_0),
.V61_1(V61_1),.V61_2(V61_2),.V61_3(V61_3),.V61_4(V61_4),.V61_5(V61_5),.V61_6(V61_6),.V61_7(V61_7),.V62_0(V62_0),.V62_1(V62_1),.V62_2(V62_2),
.V62_3(V62_3),.V62_4(V62_4),.V62_5(V62_5),.V62_6(V62_6),.V62_7(V62_7),.V63_0(V63_0),.V63_1(V63_1),.V63_2(V63_2),.V63_3(V63_3),.V63_4(V63_4),.V63_5(V63_5),.V63_6(V63_6),.V63_7(V63_7),.V64_0(V64_0),.V64_1(V64_1),.V64_2(V64_2),.V64_3(V64_3),.V64_4(V64_4),.V64_5(V64_5),.V64_6(V64_6),.V64_7(V64_7),      
      .clk(clk),.reset(reset),.prgm_b(prgm_b),.CLB_prgm_b(CLB_prgm_b),.cb_prgm_b(cb_prgm_b),.sb_prgm_b(sb_prgm_b),.io_prgm_b(io_prgm_b),.bit_in_CLB(bit_in_CLB),.bit_in_CB(bit_in_B),.bit_in_SB(bit_in_SB),.bit_in_IO(bit_in_IO),.GWE(GWE),.cb_prgm_b_in(cb_prgm_b_in),.cb_prgm_b_out(cb_prgm_b_out),.sb_prgm_b_in(sb_prgm_b_in),.sb_prgm_b_out(sb_prgm_b_out),.CLB_prgm_b_in(CLB_prgm_b_in),.CLB_prgm_b_out(CLB_prgm_b_out),.io_prgm_b_in(io_prgm_b_in),.io_prgm_b_out(io_prgm_b_out));


//For all bit-streams the bits are arranged in the decreasing order of their coordinate positions. eg. The bits belonging to the first CLB CLB_00 will be placed at the end of the CLB bitstream

initial begin

//input_file=$fopen("/home/krishna/Downloads/DEV_Git/conf_bit_stream.txt","r");
 clk = 1'b0;
 reset=1'b0; 
 prgm_b=1'b1; //indicates start of bit_stream----active low
 
 cb_prgm_b=1'b0;
 CLB_prgm_b=1'b0;
 sb_prgm_b=1'b0;
 io_prgm_b=1'b0;
 
 cb_prgm_b_in=1'b0; 
 sb_prgm_b_in=1'b0;
 CLB_prgm_b_in=1'b0;
 io_prgm_b_in=1'b0;
 
 GWE=1'b0;

 fork
/*
 #1 while(!$feof(input_file))
	begin
	CB_config_stream_final=$fscanf(input_file,"%b\n",CB_config_stream);
	SB_config_stream_final=$fscanf(input_file,"%b\n",SB_config_stream);
	CLB_config_stream_final=$fscanf(input_file,"%b\n",CLB_config_stream);
	IO_config_stream_final=$fscanf(input_file,"%b\n",IO_config_stream);
	end
	$fclose(input_file);
*/


 #1 reset=1'b1;
 #1 prgm_b=1'b0;
 
 #1 cb_prgm_b=1'b1;
 #1 cb_prgm_b_in=1'b1;
 
 #1 sb_prgm_b=1'b1;
 #1 sb_prgm_b_in=1'b1;
 
 #1 CLB_prgm_b=1'b1;
 #1 CLB_prgm_b_in=1'b1;
 
 #1 io_prgm_b_in=1'b1;
 #1 io_prgm_b=1'b1;

 #1 CB_counter=0;CB_count=0;
 #1 CLB_counter=0;CLB_count=0;
 #1 SB_counter=0;SB_count=0;
 #1 IO_counter=0;IO_count=0;
 #1 reset=1'b1;
 #2 reset=1'b0;

 join
end

initial begin
//for(i=0;i<=6074;i++)
//begin

forever #5 clk=!clk;

end

initial
begin



CB_config_stream[5119:0]= 5120'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000001000000000000000000000001000000000010000000000100000000001000000000000000000000000000000000000000000000010000000000100000000001000000000010000000000100000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000100000000000000000000000000100000000001000000000010000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001000000000010000000000000000000000000000000000000000000000000000000001000000000010000000000100000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


SB_config_stream0[7679:0]= 7680'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


SB_config_stream1[7679:0]= 7680'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


SB_config_stream2[3839:0]= 3840'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000010000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000010000000000000000000000000000000001000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



CLB_config_stream[7423:0]= 7424'b00000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000101100101000100100100000000000000001101110110000000000000010110010100010010010000000000000000110110011000000000000001011001010001001001000000000000000011011010100000000000000101100101000100100100000000000000001101110100000000000000000000000000000000000000000000001110110110000000000000000000000000000000000000000000000000110011011000000000000000000000000000000000000000000000000000101101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000101000100000011001010000000000000000101000110001000100001110101110100111100000000000000000010010101111000100010000111000111000001010000100000000000001001010111100010001000000011000100000001001010000000000000000101000110001000100000001100001100010100000000000000000010010100011000100010000000010001000000110000100000000000000001010111100010001000000011000000000001000010000000000000000101011110001000100000000100000100000000000000000000000001101110010000000010010000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000001000001000001100001100000000000001101110010000000010010000100000010000000000110000000000000001010001100010001000000010000010000001000000000000000000100101011110001000100000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000000000000000000000000000000000000000011011000000000000000000000000000000000000000000000000000001101100000000000000000000000000000000000000000000000000000110110000000000000000;

IO_config_stream[319:0]=320'b00000000000000000000000000000000000000000000000011111111000000001111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;


for(l=0;l<5120;l=l+1)
CB_config_stream_final[l]=CB_config_stream[l];

for(k=0;k<7424;k=k+1)
CLB_config_stream_final[k]=CLB_config_stream[k];


for(i0=0;i0<7680;i0=i0+1)
SB_config_stream_final[i0]=SB_config_stream0[i0];

for(i1=0;i1<7680;i1=i1+1)
SB_config_stream_final[i1+7680]=SB_config_stream1[i1];

for(i2=0;i2<3840;i2=i2+1)
SB_config_stream_final[i2+15360]=SB_config_stream2[i2];


for(m=0;m<320;m=m+1)
IO_config_stream_final[m]=IO_config_stream[m];



end

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && cb_prgm_b!=1'b0) begin
	
	
    if((CB_counter == 81) && cb_prgm_b!=1'b0) //(no of bits required for one CB) + 1= 48+1=49
	begin
	    
		CB_count=CB_count+1;
		
		CB_counter=0;
		if(CB_count==64)
		begin
			
			cb_prgm_b=1'b0;
           // prgm_b=1'b1;
			
		end
	end 
	bit_in_CB <= CB_config_stream_final[0];
	CB_config_stream_final <=CB_config_stream_final>>1;
	CB_counter=CB_counter+1;//if endsj
end 

end //always block ends


always@(posedge clk or posedge reset)
begin 

	if(prgm_b!=1'b1 && sb_prgm_b!=1'b0) begin
	
		if((SB_counter == 769) && sb_prgm_b!=1'b0) //(no of bits required for one SB +1 = 769)
			begin
	    
			SB_count=SB_count+1;
			SB_counter=0;
			if(SB_count==25)
			begin
			
				sb_prgm_b=1'b0;
		
			 prgm_b=1'b1;
			
			end
		end 
	bit_in_SB <= SB_config_stream_final[0];
	SB_config_stream_final <=SB_config_stream_final>>1;
	SB_counter=SB_counter+1;//if endsj
	end 

end //always block ends

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && CLB_prgm_b!=1'b0) 
begin

    if((CLB_counter == 465) && CLB_prgm_b!=1'b0) //(no of bits required for one CLB) + 1= 38+1=39  or (38 + (number of LUT -1))
	begin
	    
		CLB_count=CLB_count+1;
		
		CLB_counter=0;
		if(CLB_count==16)
		begin
			
			CLB_prgm_b=1'b0;
          
			
		end
	end 
	bit_in_CLB <= CLB_config_stream_final[0];
	CLB_config_stream_final <=CLB_config_stream_final>>1;
	CLB_counter=CLB_counter+1;//if endsj
end 

end //always block ends

always@(posedge clk or posedge reset)
begin 

if(prgm_b!=1'b1 && io_prgm_b!=1'b0) 
begin	
	
    if((IO_counter == 16) && io_prgm_b!=1'b0) //(no of bits required for one IO block configuration + 1= 16+1=17
	begin
	    
		IO_count=IO_count+1;
		
		IO_counter=0;
		if(IO_count==20)
		begin
			
			io_prgm_b=1'b0;
           // prgm_b=1'b1;
			
		end
	end 
	bit_in_IO <= IO_config_stream_final[0];
	IO_config_stream_final <=IO_config_stream_final>>1;
	IO_counter=IO_counter+1;//if endsj
end 

end //always block ends

//end  




initial
	begin 
#600;               //time=5 seconds
V600=1;V601=1;V602=1;V603=1;V604=1;V605=1;V606=1;V607=1;

#800;
	
V600=1;V601=1;V602=1;V603=1;V604=1;V605=1;V606=1;V607=1;

#800;
	
V600=1;V601=1;V602=1;V603=1;V604=1;V605=1;V606=1;V607=1;

#20000 $finish;
end
initial begin

    $dumpfile("test.vcd");
    $dumpvars(0,FPGA_testbench);
    $timeformat(-9, 1, " ns", 6);
	$monitor("At prgm_b=%b reset=%b SB_count=%d",prgm_b,reset,SB_count);

end

//Stimulus

endmodule
