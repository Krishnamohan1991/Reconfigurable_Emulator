`define behavioral
module switch_block(bit_in,clk,reset,prgm_b,sb_prgm_b,sb_prgm_b_in,sb_prgm_b_out,sb_prgm_b_out,A0,A1,A2,A3,A4,A5,A6,A7,B0,B1,B2,B3,B4,B5,B6,B7,
	C0,C1,C2,C3,C4,C5,C6,C7,D0,D1,D2,D3,D4,D5,D6,D7);

inout A0,A1,A2,A3,A4,A5,A6,A7,B0,B1,B2,B3,B4,B5,B6,B7,C0,C1,C2,C3,C4,C5,C6,C7,D0,D1,D2,D3,D4,D5,D6,D7;

output sb_prgm_b_out;

input bit_in,prgm_b,sb_prgm_b,sb_prgm_b_in,clk,reset;

`ifdef behavioral
 wire [1:0]A0_B0; wire [1:0]A0_B1; wire [1:0]A0_B2; wire [1:0]A0_B3; wire [1:0]A0_B4; wire [1:0]A0_B5; wire [1:0]A0_B6; wire [1:0]A0_B7; wire [1:0]A0_C0; wire [1:0]A0_C1; wire [1:0]A0_C2; wire [1:0]A0_C3; wire [1:0]A0_C4; wire [1:0]A0_C5; wire [1:0]A0_C6; wire [1:0]A0_C7; wire [1:0]A0_D0; wire [1:0]A0_D1; wire [1:0]A0_D2;wire [1:0]A0_D3; wire [1:0]A0_D4; wire [1:0]A0_D5; wire [1:0]A0_D6; wire [1:0]A0_D7; wire [1:0]A1_B0;
 wire [1:0]A1_B1; wire [1:0]A1_B2; wire [1:0]A1_B3; wire [1:0]A1_B4; wire [1:0]A1_B5; wire [1:0]A1_B6; wire [1:0]A1_B7; wire [1:0]A1_C0; wire [1:0]A1_C1; wire [1:0]A1_C2; wire [1:0]A1_C3; wire [1:0]A1_C4; wire [1:0]A1_C5; wire [1:0]A1_C6; wire [1:0]A1_C7; wire [1:0]A1_D0; wire [1:0]A1_D1; wire [1:0]A1_D2; wire [1:0]A1_D3; wire [1:0]A1_D4; wire [1:0]A1_D5; wire [1:0]A1_D6; wire [1:0]A1_D7; wire [1:0]A2_B0; wire [1:0]A2_B1;
 wire [1:0]A2_B2; wire [1:0]A2_B3; wire [1:0]A2_B4; wire [1:0]A2_B5; wire [1:0]A2_B6; wire [1:0]A2_B7; wire [1:0]A2_C0; wire [1:0]A2_C1; wire [1:0]A2_C2; wire [1:0]A2_C3; wire [1:0]A2_C4; wire [1:0]A2_C5; wire [1:0]A2_C6; wire [1:0]A2_C7; wire [1:0]A2_D0; wire [1:0]A2_D1; wire [1:0]A2_D2; wire [1:0]A2_D3; wire [1:0]A2_D4; wire [1:0]A2_D5; wire [1:0]A2_D6; wire [1:0]A2_D7; wire [1:0]A3_B0; wire [1:0]A3_B1; wire [1:0]A3_B2;
 wire [1:0]A3_B3; wire [1:0]A3_B4; wire [1:0]A3_B5; wire [1:0]A3_B6; wire [1:0]A3_B7; wire [1:0]A3_C0; wire [1:0]A3_C1; wire [1:0]A3_C2; wire [1:0]A3_C3; wire [1:0]A3_C4; wire [1:0]A3_C5; wire [1:0]A3_C6; wire [1:0]A3_C7; wire [1:0]A3_D0; wire [1:0]A3_D1; wire [1:0]A3_D2; wire [1:0]A3_D3; wire [1:0]A3_D4; wire [1:0]A3_D5; wire [1:0]A3_D6; wire [1:0]A3_D7; wire [1:0]A4_B0; wire [1:0]A4_B1; wire [1:0]A4_B2; wire [1:0]A4_B3;
 wire [1:0]A4_B4; wire [1:0]A4_B5; wire [1:0]A4_B6; wire [1:0]A4_B7; wire [1:0]A4_C0; wire [1:0]A4_C1; wire [1:0]A4_C2; wire [1:0]A4_C3; wire [1:0]A4_C4; wire [1:0]A4_C5; wire [1:0]A4_C6; wire [1:0]A4_C7; wire [1:0]A4_D0; wire [1:0]A4_D1; wire [1:0]A4_D2; wire [1:0]A4_D3; wire [1:0]A4_D4; wire [1:0]A4_D5; wire [1:0]A4_D6; wire [1:0]A4_D7; wire [1:0]A5_B0; wire [1:0]A5_B1; wire [1:0]A5_B2; wire [1:0]A5_B3; wire [1:0]A5_B4;
 wire [1:0]A5_B5; wire [1:0]A5_B6; wire [1:0]A5_B7; wire [1:0]A5_C0; wire [1:0]A5_C1; wire [1:0]A5_C2; wire [1:0]A5_C3; wire [1:0]A5_C4; wire [1:0]A5_C5; wire [1:0]A5_C6; wire [1:0]A5_C7; wire [1:0]A5_D0; wire [1:0]A5_D1; wire [1:0]A5_D2; wire [1:0]A5_D3; wire [1:0]A5_D4; wire [1:0]A5_D5; wire [1:0]A5_D6; wire [1:0]A5_D7; wire [1:0]A6_B0; wire [1:0]A6_B1; wire [1:0]A6_B2; wire [1:0]A6_B3; wire [1:0]A6_B4; wire [1:0]A6_B5;
 wire [1:0]A6_B6; wire [1:0]A6_B7; wire [1:0]A6_C0; wire [1:0]A6_C1; wire [1:0]A6_C2; wire [1:0]A6_C3; wire [1:0]A6_C4; wire [1:0]A6_C5; wire [1:0]A6_C6; wire [1:0]A6_C7; wire [1:0]A6_D0; wire [1:0]A6_D1; wire [1:0]A6_D2; wire [1:0]A6_D3; wire [1:0]A6_D4; wire [1:0]A6_D5; wire [1:0]A6_D6; wire [1:0]A6_D7; wire [1:0]A7_B0; wire [1:0]A7_B1; wire [1:0]A7_B2; wire [1:0]A7_B3; wire [1:0]A7_B4; wire [1:0]A7_B5; wire [1:0]A7_B6;
 wire [1:0]A7_B7; wire [1:0]A7_C0; wire [1:0]A7_C1; wire [1:0]A7_C2; wire [1:0]A7_C3; wire [1:0]A7_C4; wire [1:0]A7_C5; wire [1:0]A7_C6; wire [1:0]A7_C7; wire [1:0]A7_D0; wire [1:0]A7_D1; wire [1:0]A7_D2; wire [1:0]A7_D3; wire [1:0]A7_D4; wire [1:0]A7_D5; wire [1:0]A7_D6; wire [1:0]A7_D7; wire [1:0]B0_D0; wire [1:0]B0_D1; wire [1:0]B0_D2; wire [1:0]B0_D3; wire [1:0]B0_D4; wire [1:0]B0_D5; wire [1:0]B0_D6; wire [1:0]B0_D7;
 wire [1:0]B0_C0; wire [1:0]B0_C1; wire [1:0]B0_C2; wire [1:0]B0_C3; wire [1:0]B0_C4; wire [1:0]B0_C5; wire [1:0]B0_C6; wire [1:0]B0_C7; wire [1:0]B1_D0; wire [1:0]B1_D1; wire [1:0]B1_D2; wire [1:0]B1_D3; wire [1:0]B1_D4; wire [1:0]B1_D5; wire [1:0]B1_D6; wire [1:0]B1_D7; wire [1:0]B1_C0; wire [1:0]B1_C1; wire [1:0]B1_C2; wire [1:0]B1_C3; wire [1:0]B1_C4; wire [1:0]B1_C5; wire [1:0]B1_C6; wire [1:0]B1_C7; wire [1:0]B2_D0;
 wire [1:0]B2_D1; wire [1:0]B2_D2; wire [1:0]B2_D3; wire [1:0]B2_D4; wire [1:0]B2_D5; wire [1:0]B2_D6; wire [1:0]B2_D7; wire [1:0]B2_C0; wire [1:0]B2_C1; wire [1:0]B2_C2; wire [1:0]B2_C3; wire [1:0]B2_C4; wire [1:0]B2_C5; wire [1:0]B2_C6; wire [1:0]B2_C7; wire [1:0]B3_D0; wire [1:0]B3_D1; wire [1:0]B3_D2; wire [1:0]B3_D3; wire [1:0]B3_D4; wire [1:0]B3_D5; wire [1:0]B3_D6; wire [1:0]B3_D7; wire [1:0]B3_C0; wire [1:0]B3_C1;
 wire [1:0]B3_C2; wire [1:0]B3_C3; wire [1:0]B3_C4; wire [1:0]B3_C5; wire [1:0]B3_C6; wire [1:0]B3_C7; wire [1:0]B4_D0; wire [1:0]B4_D1; wire [1:0]B4_D2; wire [1:0]B4_D3; wire [1:0]B4_D4; wire [1:0]B4_D5; wire [1:0]B4_D6; wire [1:0]B4_D7; wire [1:0]B4_C0; wire [1:0]B4_C1; wire [1:0]B4_C2; wire [1:0]B4_C3; wire [1:0]B4_C4; wire [1:0]B4_C5; wire [1:0]B4_C6; wire [1:0]B4_C7; wire [1:0]B5_D0; wire [1:0]B5_D1; wire [1:0]B5_D2;
 wire [1:0]B5_D3; wire [1:0]B5_D4; wire [1:0]B5_D5; wire [1:0]B5_D6; wire [1:0]B5_D7; wire [1:0]B5_C0; wire [1:0]B5_C1; wire [1:0]B5_C2; wire [1:0]B5_C3; wire [1:0]B5_C4; wire [1:0]B5_C5; wire [1:0]B5_C6; wire [1:0]B5_C7; wire [1:0]B6_D0; wire [1:0]B6_D1; wire [1:0]B6_D2; wire [1:0]B6_D3; wire [1:0]B6_D4; wire [1:0]B6_D5; wire [1:0]B6_D6; wire [1:0]B6_D7; wire [1:0]B6_C0; wire [1:0]B6_C1; wire [1:0]B6_C2; wire [1:0]B6_C3;
 wire [1:0]B6_C4; wire [1:0]B6_C5; wire [1:0]B6_C6; wire [1:0]B6_C7; wire [1:0]B7_D0; wire [1:0]B7_D1; wire [1:0]B7_D2; wire [1:0]B7_D3; wire [1:0]B7_D4; wire [1:0]B7_D5; wire [1:0]B7_D6; wire [1:0]B7_D7; wire [1:0]B7_C0; wire [1:0]B7_C1; wire [1:0]B7_C2; wire [1:0]B7_C3; wire [1:0]B7_C4; wire [1:0]B7_C5; wire [1:0]B7_C6; wire [1:0]B7_C7; wire [1:0]C0_D0; wire [1:0]C0_D1; wire [1:0]C0_D2; wire [1:0]C0_D3; wire [1:0]C0_D4;
 wire [1:0]C0_D5; wire [1:0]C0_D6; wire [1:0]C0_D7; wire [1:0]C1_D0; wire [1:0]C1_D1; wire [1:0]C1_D2; wire [1:0]C1_D3; wire [1:0]C1_D4; wire [1:0]C1_D5; wire [1:0]C1_D6; wire [1:0]C1_D7; wire [1:0]C2_D0; wire [1:0]C2_D1; wire [1:0]C2_D2; wire [1:0]C2_D3; wire [1:0]C2_D4; wire [1:0]C2_D5; wire [1:0]C2_D6; wire [1:0]C2_D7; wire [1:0]C3_D0; wire [1:0]C3_D1; wire [1:0]C3_D2; wire [1:0]C3_D3; wire [1:0]C3_D4; wire [1:0]C3_D5;
 wire [1:0]C3_D6; wire [1:0]C3_D7; wire [1:0]C4_D0; wire [1:0]C4_D1; wire [1:0]C4_D2; wire [1:0]C4_D3; wire [1:0]C4_D4; wire [1:0]C4_D5; wire [1:0]C4_D6; wire [1:0]C4_D7; wire [1:0]C5_D0; wire [1:0]C5_D1; wire [1:0]C5_D2; wire [1:0]C5_D3; wire [1:0]C5_D4; wire [1:0]C5_D5; wire [1:0]C5_D6; wire [1:0]C5_D7; wire [1:0]C6_D0; wire [1:0]C6_D1; wire [1:0]C6_D2; wire [1:0]C6_D3; wire [1:0]C6_D4; wire [1:0]C6_D5; wire [1:0]C6_D6;
 wire [1:0]C6_D7; wire [1:0]C7_D0; wire [1:0]C7_D1; wire [1:0]C7_D2; wire [1:0]C7_D3; wire [1:0]C7_D4; wire [1:0]C7_D5; wire [1:0]C7_D6; wire [1:0]C7_D7;


SB_config_behav SB_behav_config(.bit_in(bit_in),.prgm_b(prgm_b),.sb_prgm_b(sb_prgm_b),.clk(clk),.reset(reset),.sb_prgm_b_in(sb_prgm_b_in),.sb_prgm_b_out(sb_prgm_b_out),
.A0_B0(A0_B0),.A0_B1(A0_B1),.A0_B2(A0_B2),.A0_B3(A0_B3),.A0_B4(A0_B4),.A0_B5(A0_B5),.A0_B6(A0_B6),.A0_B7(A0_B7),.A0_C0(A0_C0),.A0_C1(A0_C1),.A0_C2(A0_C2),.A0_C3(A0_C3),.A0_C4(A0_C4),.A0_C5(A0_C5),.A0_C6(A0_C6),.A0_C7(A0_C7),.A0_D0(A0_D0),.A0_D1(A0_D1),.A0_D2(A0_D2),.A0_D3(A0_D3),.A0_D4(A0_D4),.A0_D5(A0_D5),.A0_D6(A0_D6),.A0_D7(A0_D7),.A1_B0(A1_B0),
.A1_B1(A1_B1),.A1_B2(A1_B2),.A1_B3(A1_B3),.A1_B4(A1_B4),.A1_B5(A1_B5),.A1_B6(A1_B6),.A1_B7(A1_B7),.A1_C0(A1_C0),.A1_C1(A1_C1),.A1_C2(A1_C2),.A1_C3(A1_C3),.A1_C4(A1_C4),.A1_C5(A1_C5),.A1_C6(A1_C6),.A1_C7(A1_C7),.A1_D0(A1_D0),.A1_D1(A1_D1),.A1_D2(A1_D2),.A1_D3(A1_D3),.A1_D4(A1_D4),.A1_D5(A1_D5),.A1_D6(A1_D6),.A1_D7(A1_D7),.A2_B0(A2_B0),.A2_B1(A2_B1),
.A2_B2(A2_B2),.A2_B3(A2_B3),.A2_B4(A2_B4),.A2_B5(A2_B5),.A2_B6(A2_B6),.A2_B7(A2_B7),.A2_C0(A2_C0),.A2_C1(A2_C1),.A2_C2(A2_C2),.A2_C3(A2_C3),.A2_C4(A2_C4),.A2_C5(A2_C5),.A2_C6(A2_C6),.A2_C7(A2_C7),.A2_D0(A2_D0),.A2_D1(A2_D1),.A2_D2(A2_D2),.A2_D3(A2_D3),.A2_D4(A2_D4),.A2_D5(A2_D5),.A2_D6(A2_D6),.A2_D7(A2_D7),.A3_B0(A3_B0),.A3_B1(A3_B1),.A3_B2(A3_B2),
.A3_B3(A3_B3),.A3_B4(A3_B4),.A3_B5(A3_B5),.A3_B6(A3_B6),.A3_B7(A3_B7),.A3_C0(A3_C0),.A3_C1(A3_C1),.A3_C2(A3_C2),.A3_C3(A3_C3),.A3_C4(A3_C4),.A3_C5(A3_C5),.A3_C6(A3_C6),.A3_C7(A3_C7),.A3_D0(A3_D0),.A3_D1(A3_D1),.A3_D2(A3_D2),.A3_D3(A3_D3),.A3_D4(A3_D4),.A3_D5(A3_D5),.A3_D6(A3_D6),.A3_D7(A3_D7),.A4_B0(A4_B0),.A4_B1(A4_B1),.A4_B2(A4_B2),.A4_B3(A4_B3),
.A4_B4(A4_B4),.A4_B5(A4_B5),.A4_B6(A4_B6),.A4_B7(A4_B7),.A4_C0(A4_C0),.A4_C1(A4_C1),.A4_C2(A4_C2),.A4_C3(A4_C3),.A4_C4(A4_C4),.A4_C5(A4_C5),.A4_C6(A4_C6),.A4_C7(A4_C7),.A4_D0(A4_D0),.A4_D1(A4_D1),.A4_D2(A4_D2),.A4_D3(A4_D3),.A4_D4(A4_D4),.A4_D5(A4_D5),.A4_D6(A4_D6),.A4_D7(A4_D7),.A5_B0(A5_B0),.A5_B1(A5_B1),.A5_B2(A5_B2),.A5_B3(A5_B3),.A5_B4(A5_B4),
.A5_B5(A5_B5),.A5_B6(A5_B6),.A5_B7(A5_B7),.A5_C0(A5_C0),.A5_C1(A5_C1),.A5_C2(A5_C2),.A5_C3(A5_C3),.A5_C4(A5_C4),.A5_C5(A5_C5),.A5_C6(A5_C6),.A5_C7(A5_C7),.A5_D0(A5_D0),.A5_D1(A5_D1),.A5_D2(A5_D2),.A5_D3(A5_D3),.A5_D4(A5_D4),.A5_D5(A5_D5),.A5_D6(A5_D6),.A5_D7(A5_D7),.A6_B0(A6_B0),.A6_B1(A6_B1),.A6_B2(A6_B2),.A6_B3(A6_B3),.A6_B4(A6_B4),.A6_B5(A6_B5),
.A6_B6(A6_B6),.A6_B7(A6_B7),.A6_C0(A6_C0),.A6_C1(A6_C1),.A6_C2(A6_C2),.A6_C3(A6_C3),.A6_C4(A6_C4),.A6_C5(A6_C5),.A6_C6(A6_C6),.A6_C7(A6_C7),.A6_D0(A6_D0),.A6_D1(A6_D1),.A6_D2(A6_D2),.A6_D3(A6_D3),.A6_D4(A6_D4),.A6_D5(A6_D5),.A6_D6(A6_D6),.A6_D7(A6_D7),.A7_B0(A7_B0),.A7_B1(A7_B1),.A7_B2(A7_B2),.A7_B3(A7_B3),.A7_B4(A7_B4),.A7_B5(A7_B5),.A7_B6(A7_B6),
.A7_B7(A7_B7),.A7_C0(A7_C0),.A7_C1(A7_C1),.A7_C2(A7_C2),.A7_C3(A7_C3),.A7_C4(A7_C4),.A7_C5(A7_C5),.A7_C6(A7_C6),.A7_C7(A7_C7),.A7_D0(A7_D0),.A7_D1(A7_D1),.A7_D2(A7_D2),.A7_D3(A7_D3),.A7_D4(A7_D4),.A7_D5(A7_D5),.A7_D6(A7_D6),.A7_D7(A7_D7),.B0_D0(B0_D0),.B0_D1(B0_D1),.B0_D2(B0_D2),.B0_D3(B0_D3),.B0_D4(B0_D4),.B0_D5(B0_D5),.B0_D6(B0_D6),.B0_D7(B0_D7),
.B0_C0(B0_C0),.B0_C1(B0_C1),.B0_C2(B0_C2),.B0_C3(B0_C3),.B0_C4(B0_C4),.B0_C5(B0_C5),.B0_C6(B0_C6),.B0_C7(B0_C7),.B1_D0(B1_D0),.B1_D1(B1_D1),.B1_D2(B1_D2),.B1_D3(B1_D3),.B1_D4(B1_D4),.B1_D5(B1_D5),.B1_D6(B1_D6),.B1_D7(B1_D7),.B1_C0(B1_C0),.B1_C1(B1_C1),.B1_C2(B1_C2),.B1_C3(B1_C3),.B1_C4(B1_C4),.B1_C5(B1_C5),.B1_C6(B1_C6),.B1_C7(B1_C7),.B2_D0(B2_D0),
.B2_D1(B2_D1),.B2_D2(B2_D2),.B2_D3(B2_D3),.B2_D4(B2_D4),.B2_D5(B2_D5),.B2_D6(B2_D6),.B2_D7(B2_D7),.B2_C0(B2_C0),.B2_C1(B2_C1),.B2_C2(B2_C2),.B2_C3(B2_C3),.B2_C4(B2_C4),.B2_C5(B2_C5),.B2_C6(B2_C6),.B2_C7(B2_C7),.B3_D0(B3_D0),.B3_D1(B3_D1),.B3_D2(B3_D2),.B3_D3(B3_D3),.B3_D4(B3_D4),.B3_D5(B3_D5),.B3_D6(B3_D6),.B3_D7(B3_D7),.B3_C0(B3_C0),.B3_C1(B3_C1),
.B3_C2(B3_C2),.B3_C3(B3_C3),.B3_C4(B3_C4),.B3_C5(B3_C5),.B3_C6(B3_C6),.B3_C7(B3_C7),.B4_D0(B4_D0),.B4_D1(B4_D1),.B4_D2(B4_D2),.B4_D3(B4_D3),.B4_D4(B4_D4),.B4_D5(B4_D5),.B4_D6(B4_D6),.B4_D7(B4_D7),.B4_C0(B4_C0),.B4_C1(B4_C1),.B4_C2(B4_C2),.B4_C3(B4_C3),.B4_C4(B4_C4),.B4_C5(B4_C5),.B4_C6(B4_C6),.B4_C7(B4_C7),.B5_D0(B5_D0),.B5_D1(B5_D1),.B5_D2(B5_D2),
.B5_D3(B5_D3),.B5_D4(B5_D4),.B5_D5(B5_D5),.B5_D6(B5_D6),.B5_D7(B5_D7),.B5_C0(B5_C0),.B5_C1(B5_C1),.B5_C2(B5_C2),.B5_C3(B5_C3),.B5_C4(B5_C4),.B5_C5(B5_C5),.B5_C6(B5_C6),.B5_C7(B5_C7),.B6_D0(B6_D0),.B6_D1(B6_D1),.B6_D2(B6_D2),.B6_D3(B6_D3),.B6_D4(B6_D4),.B6_D5(B6_D5),.B6_D6(B6_D6),.B6_D7(B6_D7),.B6_C0(B6_C0),.B6_C1(B6_C1),.B6_C2(B6_C2),.B6_C3(B6_C3),
.B6_C4(B6_C4),.B6_C5(B6_C5),.B6_C6(B6_C6),.B6_C7(B6_C7),.B7_D0(B7_D0),.B7_D1(B7_D1),.B7_D2(B7_D2),.B7_D3(B7_D3),.B7_D4(B7_D4),.B7_D5(B7_D5),.B7_D6(B7_D6),.B7_D7(B7_D7),.B7_C0(B7_C0),.B7_C1(B7_C1),.B7_C2(B7_C2),.B7_C3(B7_C3),.B7_C4(B7_C4),.B7_C5(B7_C5),.B7_C6(B7_C6),.B7_C7(B7_C7),.C0_D0(C0_D0),.C0_D1(C0_D1),.C0_D2(C0_D2),.C0_D3(C0_D3),.C0_D4(C0_D4),
.C0_D5(C0_D5),.C0_D6(C0_D6),.C0_D7(C0_D7),.C1_D0(C1_D0),.C1_D1(C1_D1),.C1_D2(C1_D2),.C1_D3(C1_D3),.C1_D4(C1_D4),.C1_D5(C1_D5),.C1_D6(C1_D6),.C1_D7(C1_D7),.C2_D0(C2_D0),.C2_D1(C2_D1),.C2_D2(C2_D2),.C2_D3(C2_D3),.C2_D4(C2_D4),.C2_D5(C2_D5),.C2_D6(C2_D6),.C2_D7(C2_D7),.C3_D0(C3_D0),.C3_D1(C3_D1),.C3_D2(C3_D2),.C3_D3(C3_D3),.C3_D4(C3_D4),.C3_D5(C3_D5),
.C3_D6(C3_D6),.C3_D7(C3_D7),.C4_D0(C4_D0),.C4_D1(C4_D1),.C4_D2(C4_D2),.C4_D3(C4_D3),.C4_D4(C4_D4),.C4_D5(C4_D5),.C4_D6(C4_D6),.C4_D7(C4_D7),.C5_D0(C5_D0),.C5_D1(C5_D1),.C5_D2(C5_D2),.C5_D3(C5_D3),.C5_D4(C5_D4),.C5_D5(C5_D5),.C5_D6(C5_D6),.C5_D7(C5_D7),.C6_D0(C6_D0),.C6_D1(C6_D1),.C6_D2(C6_D2),.C6_D3(C6_D3),.C6_D4(C6_D4),.C6_D5(C6_D5),.C6_D6(C6_D6),
.C6_D7(C6_D7),.C7_D0(C7_D0),.C7_D1(C7_D1),.C7_D2(C7_D2),.C7_D3(C7_D3),.C7_D4(C7_D4),.C7_D5(C7_D5),.C7_D6(C7_D6),.C7_D7(C7_D7));




bidir_switch A0B0(.port1(A0),.port2(B0),.enable_dir(A0_B0));    bidir_switch A1B0(.port1(A1),.port2(B0),.enable_dir(A1_B0));  bidir_switch SC1(.port1(A2),.port2(B0),.enable_dir(A2_B0));   bidir_switch SD1(.port1(A3),.port2(B0),.enable_dir(A3_B0));
                                                                              
bidir_switch A0B1(.port1(A0),.port2(B1),.enable_dir(A0_B1));    bidir_switch A1B1(.port1(A1),.port2(B1),.enable_dir(A1_B1));   bidir_switch SC2(.port1(A2),.port2(B1),.enable_dir(A2_B1));   bidir_switch SD2(.port1(A3),.port2(B1),.enable_dir(A3_B1));
                                                                              
bidir_switch A0B2(.port1(A0),.port2(B2),.enable_dir(A0_B2));    bidir_switch A1B2(.port1(A1),.port2(B2),.enable_dir(A1_B2));   bidir_switch SC3(.port1(A2),.port2(B2),.enable_dir(A2_B2));   bidir_switch SD3(.port1(A3),.port2(B2),.enable_dir(A3_B2));
                                                                              
bidir_switch A0B3(.port1(A0),.port2(B3),.enable_dir(A0_B3));    bidir_switch A1B3(.port1(A1),.port2(B3),.enable_dir(A1_B3));   bidir_switch SC4(.port1(A2),.port2(B3),.enable_dir(A2_B3));   bidir_switch SD4(.port1(A3),.port2(B3),.enable_dir(A3_B3));
                                                                              
bidir_switch A0B4(.port1(A0),.port2(B4),.enable_dir(A0_B4));    bidir_switch A1B4(.port1(A1),.port2(B4),.enable_dir(A1_B4));   bidir_switch SC5(.port1(A2),.port2(B4),.enable_dir(A2_B4));   bidir_switch SD5(.port1(A3),.port2(B4),.enable_dir(A3_B4));
                                                                              
bidir_switch A0B5(.port1(A0),.port2(B5),.enable_dir(A0_B5));    bidir_switch A1B5(.port1(A1),.port2(B5),.enable_dir(A1_B5));   bidir_switch SC6(.port1(A2),.port2(B5),.enable_dir(A2_B5));   bidir_switch SD6(.port1(A3),.port2(B5),.enable_dir(A3_B5));
                                                                              
bidir_switch A0B6(.port1(A0),.port2(B6),.enable_dir(A0_B6));    bidir_switch A1B6(.port1(A1),.port2(B6),.enable_dir(A1_B6));   bidir_switch SC7(.port1(A2),.port2(B6),.enable_dir(A2_B6));   bidir_switch SD7(.port1(A3),.port2(B6),.enable_dir(A3_B6));
                                                                              
bidir_switch A0B7(.port1(A0),.port2(B7),.enable_dir(A0_B7));    bidir_switch A1B7(.port1(A1),.port2(B7),.enable_dir(A1_B7));   bidir_switch SC8(.port1(A2),.port2(B7),.enable_dir(A2_B7));   bidir_switch SD8(.port1(A3),.port2(B7),.enable_dir(A3_B7));
              
bidir_switch A0C0(.port1(A0),.port2(C0),.enable_dir(A0_C0));   bidir_switch A1C0(.port1(A1),.port2(C0),.enable_dir(A1_C0));   bidir_switch SC9(.port1(A2),.port2(C0),.enable_dir(A2_C0));   bidir_switch SD9(.port1(A3),.port2(C0),.enable_dir(A3_C0));
                                                                             
bidir_switch A0C1(.port1(A0),.port2(C1),.enable_dir(A0_C1));   bidir_switch A1C1(.port1(A1),.port2(C1),.enable_dir(A1_C1));  bidir_switch SC10(.port1(A2),.port2(C1),.enable_dir(A2_C1));  bidir_switch SD10(.port1(A3),.port2(C1),.enable_dir(A3_C1));
                                                                             
bidir_switch A0C2(.port1(A0),.port2(C2),.enable_dir(A0_C2));   bidir_switch A1C2(.port1(A1),.port2(C2),.enable_dir(A1_C2));  bidir_switch SC11(.port1(A2),.port2(C2),.enable_dir(A2_C2));  bidir_switch SD11(.port1(A3),.port2(C2),.enable_dir(A3_C2));
                                                                             
bidir_switch A0C3(.port1(A0),.port2(C3),.enable_dir(A0_C3));   bidir_switch A1C3(.port1(A1),.port2(C3),.enable_dir(A1_C3));  bidir_switch SC12(.port1(A2),.port2(C3),.enable_dir(A2_C3));  bidir_switch SD12(.port1(A3),.port2(C3),.enable_dir(A3_C3));
                                                                             
bidir_switch A0C4(.port1(A0),.port2(C4),.enable_dir(A0_C4));   bidir_switch A1C4(.port1(A1),.port2(C4),.enable_dir(A1_C4));  bidir_switch SC13(.port1(A2),.port2(C4),.enable_dir(A2_C4));  bidir_switch SD13(.port1(A3),.port2(C4),.enable_dir(A3_C4));
                                                                             
bidir_switch A0C5(.port1(A0),.port2(C5),.enable_dir(A0_C5));   bidir_switch A1C5(.port1(A1),.port2(C5),.enable_dir(A1_C5));  bidir_switch SC14(.port1(A2),.port2(C5),.enable_dir(A2_C5));  bidir_switch SD14(.port1(A3),.port2(C5),.enable_dir(A3_C5));
                                                                             
bidir_switch A0C6(.port1(A0),.port2(C6),.enable_dir(A0_C6));   bidir_switch A1C6(.port1(A1),.port2(C6),.enable_dir(A1_C6));  bidir_switch SC15(.port1(A2),.port2(C6),.enable_dir(A2_C6));  bidir_switch SD15(.port1(A3),.port2(C6),.enable_dir(A3_C6));
                                                                             
bidir_switch A0C7(.port1(A0),.port2(C7),.enable_dir(A0_C7));   bidir_switch A1C7(.port1(A1),.port2(C7),.enable_dir(A1_C7));  bidir_switch SC16(.port1(A2),.port2(C7),.enable_dir(A2_C7));  bidir_switch SD16(.port1(A3),.port2(C7),.enable_dir(A3_C7));
              
bidir_switch A0D0(.port1(A0),.port2(D0),.enable_dir(A0_D0));   bidir_switch A1D0(.port1(A1),.port2(D0),.enable_dir(A1_D0));  bidir_switch SC17(.port1(A2),.port2(D0),.enable_dir(A2_D0));  bidir_switch SD17(.port1(A3),.port2(D0),.enable_dir(A3_D0));
              
bidir_switch A0D1(.port1(A0),.port2(D1),.enable_dir(A0_D1));   bidir_switch A1D1(.port1(A1),.port2(D1),.enable_dir(A1_D1));  bidir_switch SC18(.port1(A2),.port2(D1),.enable_dir(A2_D1));  bidir_switch SD18(.port1(A3),.port2(D1),.enable_dir(A3_D1));
                                                                              
bidir_switch A0D2(.port1(A0),.port2(D2),.enable_dir(A0_D2));   bidir_switch A1D2(.port1(A1),.port2(D2),.enable_dir(A1_D2));  bidir_switch SC19(.port1(A2),.port2(D2),.enable_dir(A2_D2));  bidir_switch SD19(.port1(A3),.port2(D2),.enable_dir(A3_D2));
                                                                              
bidir_switch A0D3(.port1(A0),.port2(D3),.enable_dir(A0_D3));   bidir_switch A1D3(.port1(A1),.port2(D3),.enable_dir(A1_D3));  bidir_switch SC20(.port1(A2),.port2(D3),.enable_dir(A2_D3));  bidir_switch SD20(.port1(A3),.port2(D3),.enable_dir(A3_D3));
                                                                              
bidir_switch A0D4(.port1(A0),.port2(D4),.enable_dir(A0_D4));   bidir_switch A1D4(.port1(A1),.port2(D4),.enable_dir(A1_D4));  bidir_switch SC21(.port1(A2),.port2(D4),.enable_dir(A2_D4));  bidir_switch SD21(.port1(A3),.port2(D4),.enable_dir(A3_D4));
                                                                              
bidir_switch A0D5(.port1(A0),.port2(D5),.enable_dir(A0_D5));   bidir_switch A1D5(.port1(A1),.port2(D5),.enable_dir(A1_D5));  bidir_switch SC22(.port1(A2),.port2(D5),.enable_dir(A2_D5));  bidir_switch SD22(.port1(A3),.port2(D5),.enable_dir(A3_D5));
                                                                              
bidir_switch A0D6(.port1(A0),.port2(D6),.enable_dir(A0_D6));   bidir_switch A1D6(.port1(A1),.port2(D6),.enable_dir(A1_D6));  bidir_switch SC23(.port1(A2),.port2(D6),.enable_dir(A2_D6));  bidir_switch SD23(.port1(A3),.port2(D6),.enable_dir(A3_D6));
                                                                              
bidir_switch A0D7(.port1(A0),.port2(D7),.enable_dir(A0_D7));   bidir_switch A1D7(.port1(A1),.port2(D7),.enable_dir(A1_D7));  bidir_switch SC24(.port1(A2),.port2(D7),.enable_dir(A2_D7));  bidir_switch SD24(.port1(A3),.port2(D7),.enable_dir(A3_D7));






bidir_switch SE1(.port1(A4),.port2(B0),.enable_dir(A4_B0));	   bidir_switch SG1(.port1(B0),.port2(A5),.enable_dir(A5_B0));   bidir_switch SH1(.port1(B0),.port2(A6),.enable_dir(A6_B0));	bidir_switch SI1(.port1(B0),.port2(A7),.enable_dir(A7_B0));

bidir_switch SE2(.port1(A4),.port2(B1),.enable_dir(A4_B1));    bidir_switch SG2(.port1(B1),.port2(A5),.enable_dir(A5_B1));   bidir_switch SH2(.port1(B1),.port2(A6),.enable_dir(A6_B1));    bidir_switch SI2(.port1(B1),.port2(A7),.enable_dir(A7_B1));

bidir_switch SE3(.port1(A4),.port2(B2),.enable_dir(A4_B2));    bidir_switch SG3(.port1(B2),.port2(A5),.enable_dir(A5_B2));   bidir_switch SH3(.port1(B2),.port2(A6),.enable_dir(A6_B2));    bidir_switch SI3(.port1(B2),.port2(A7),.enable_dir(A7_B2));

bidir_switch SE4(.port1(A4),.port2(B3),.enable_dir(A4_B3));    bidir_switch SG4(.port1(B3),.port2(A5),.enable_dir(A5_B3));   bidir_switch SH4(.port1(B3),.port2(A6),.enable_dir(A6_B3));    bidir_switch SI4(.port1(B3),.port2(A7),.enable_dir(A7_B3));

bidir_switch SE5(.port1(A4),.port2(B4),.enable_dir(A4_B4));    bidir_switch SG5(.port1(B4),.port2(A5),.enable_dir(A5_B4));   bidir_switch SH5(.port1(B4),.port2(A6),.enable_dir(A6_B4));    bidir_switch SI5(.port1(B4),.port2(A7),.enable_dir(A7_B4));

bidir_switch SE6(.port1(A4),.port2(B5),.enable_dir(A4_B5));    bidir_switch SG6(.port1(B5),.port2(A5),.enable_dir(A5_B5));   bidir_switch SH6(.port1(B5),.port2(A6),.enable_dir(A6_B5));    bidir_switch SI6(.port1(B5),.port2(A7),.enable_dir(A7_B5));

bidir_switch SE7(.port1(A4),.port2(B6),.enable_dir(A4_B6));    bidir_switch SG7(.port1(B6),.port2(A5),.enable_dir(A5_B6));   bidir_switch SH7(.port1(B6),.port2(A6),.enable_dir(A6_B6));    bidir_switch SI7(.port1(B6),.port2(A7),.enable_dir(A7_B6));

bidir_switch SE8(.port1(A4),.port2(B7),.enable_dir(A4_B7));    bidir_switch SG8(.port1(B7),.port2(A5),.enable_dir(A5_B7));   bidir_switch SH8(.port1(B7),.port2(A6),.enable_dir(A6_B7));    bidir_switch SI8(.port1(B7),.port2(A7),.enable_dir(A7_B7));

bidir_switch SE9(.port1(A4),.port2(C0),.enable_dir(A4_C0));    bidir_switch SG9(.port1(C0),.port2(A5),.enable_dir(A5_C0));   bidir_switch SH9(.port1(C0),.port2(A6),.enable_dir(A6_C0));    bidir_switch SI9(.port1(C0),.port2(A7),.enable_dir(A7_C0));

bidir_switch SE10(.port1(A4),.port2(C1),.enable_dir(A4_C1));   bidir_switch SG10(.port1(C1),.port2(A5),.enable_dir(A5_C1));  bidir_switch SH10(.port1(C1),.port2(A6),.enable_dir(A6_C1));   bidir_switch SI10(.port1(C1),.port2(A7),.enable_dir(A7_C1));

bidir_switch SE11(.port1(A4),.port2(C2),.enable_dir(A4_C2));   bidir_switch SG11(.port1(C2),.port2(A5),.enable_dir(A5_C2));  bidir_switch SH11(.port1(C2),.port2(A6),.enable_dir(A6_C2));   bidir_switch SI11(.port1(C2),.port2(A7),.enable_dir(A7_C2));

bidir_switch SE12(.port1(A4),.port2(C3),.enable_dir(A4_C3));   bidir_switch SG12(.port1(C3),.port2(A5),.enable_dir(A5_C3));  bidir_switch SH12(.port1(C3),.port2(A6),.enable_dir(A6_C3));   bidir_switch SI12(.port1(C3),.port2(A7),.enable_dir(A7_C3));

bidir_switch SE13(.port1(A4),.port2(C4),.enable_dir(A4_C4));   bidir_switch SG13(.port1(C4),.port2(A5),.enable_dir(A5_C4));  bidir_switch SH13(.port1(C4),.port2(A6),.enable_dir(A6_C4));   bidir_switch SI13(.port1(C4),.port2(A7),.enable_dir(A7_C4));

bidir_switch SE14(.port1(A4),.port2(C5),.enable_dir(A4_C5));   bidir_switch SG14(.port1(C5),.port2(A5),.enable_dir(A5_C5));  bidir_switch SH14(.port1(C5),.port2(A6),.enable_dir(A6_C5));   bidir_switch SI14(.port1(C5),.port2(A7),.enable_dir(A7_C5));

bidir_switch SE15(.port1(A4),.port2(C6),.enable_dir(A4_C6));   bidir_switch SG15(.port1(C6),.port2(A5),.enable_dir(A5_C6));  bidir_switch SH15(.port1(C6),.port2(A6),.enable_dir(A6_C6));   bidir_switch SI15(.port1(C6),.port2(A7),.enable_dir(A7_C6));

bidir_switch SE16(.port1(A4),.port2(C7),.enable_dir(A4_C7));   bidir_switch SG16(.port1(C7),.port2(A5),.enable_dir(A5_C7));  bidir_switch SH16(.port1(C7),.port2(A6),.enable_dir(A6_C7));   bidir_switch SI16(.port1(C7),.port2(A7),.enable_dir(A7_C7));

bidir_switch SE17(.port1(A4),.port2(D0),.enable_dir(A4_D0));   bidir_switch SG17(.port1(D0),.port2(A5),.enable_dir(A5_D0));  bidir_switch SH17(.port1(D0),.port2(A6),.enable_dir(A6_D0));   bidir_switch SI17(.port1(D0),.port2(A7),.enable_dir(A7_D0));

bidir_switch SE18(.port1(A4),.port2(D1),.enable_dir(A4_D1));   bidir_switch SG18(.port1(D1),.port2(A5),.enable_dir(A5_D1));  bidir_switch SH18(.port1(D1),.port2(A6),.enable_dir(A6_D1));   bidir_switch SI18(.port1(D1),.port2(A7),.enable_dir(A7_D1));

bidir_switch SE19(.port1(A4),.port2(D2),.enable_dir(A4_D2));   bidir_switch SG19(.port1(D2),.port2(A5),.enable_dir(A5_D2));  bidir_switch SH19(.port1(D2),.port2(A6),.enable_dir(A6_D2));   bidir_switch SI19(.port1(D2),.port2(A7),.enable_dir(A7_D2));

bidir_switch SE20(.port1(A4),.port2(D3),.enable_dir(A4_D3));   bidir_switch SG20(.port1(D3),.port2(A5),.enable_dir(A5_D3));  bidir_switch SH20(.port1(D3),.port2(A6),.enable_dir(A6_D3));   bidir_switch SI20(.port1(D3),.port2(A7),.enable_dir(A7_D3));

bidir_switch SE21(.port1(A4),.port2(D4),.enable_dir(A4_D4));   bidir_switch SG21(.port1(D4),.port2(A5),.enable_dir(A5_D4));  bidir_switch SH21(.port1(D4),.port2(A6),.enable_dir(A6_D4));   bidir_switch SI21(.port1(D4),.port2(A7),.enable_dir(A7_D4));

bidir_switch SE22(.port1(A4),.port2(D5),.enable_dir(A4_D5));   bidir_switch SG22(.port1(D5),.port2(A5),.enable_dir(A5_D5));  bidir_switch SH22(.port1(D5),.port2(A6),.enable_dir(A6_D5));   bidir_switch SI22(.port1(D5),.port2(A7),.enable_dir(A7_D5));

bidir_switch SE23(.port1(A4),.port2(D6),.enable_dir(A4_D6));   bidir_switch SG23(.port1(D6),.port2(A5),.enable_dir(A5_D6));  bidir_switch SH23(.port1(D6),.port2(A6),.enable_dir(A6_D6));   bidir_switch SI23(.port1(D6),.port2(A7),.enable_dir(A7_D6));

bidir_switch SE24(.port1(A4),.port2(D7),.enable_dir(A4_D7));   bidir_switch SG24(.port1(D7),.port2(A5),.enable_dir(A5_D7));  bidir_switch SH24(.port1(D7),.port2(A6),.enable_dir(A6_D7));   bidir_switch SI24(.port1(D7),.port2(A7),.enable_dir(A7_D7));

             

             

bidir_switch SJ1(.port1(B0),.port2(D0),.enable_dir(B0_D0));	  bidir_switch SK1(.port1(B1),.port2(D0),.enable_dir(B1_D0));   bidir_switch SL1(.port1(B2),.port2(D0),.enable_dir(B2_D0));   bidir_switch SM1(.port1(B3),.port2(D0),.enable_dir(B3_D0));

bidir_switch SJ2(.port1(B0),.port2(D1),.enable_dir(B0_D1));   bidir_switch SK2(.port1(B1),.port2(D1),.enable_dir(B1_D1));   bidir_switch SL2(.port1(B2),.port2(D1),.enable_dir(B2_D1));   bidir_switch SM2(.port1(B3),.port2(D1),.enable_dir(B3_D1));

bidir_switch SJ3(.port1(B0),.port2(D2),.enable_dir(B0_D2));   bidir_switch SK3(.port1(B1),.port2(D2),.enable_dir(B1_D2));   bidir_switch SL3(.port1(B2),.port2(D2),.enable_dir(B2_D2));   bidir_switch SM3(.port1(B3),.port2(D2),.enable_dir(B3_D2));

bidir_switch SJ4(.port1(B0),.port2(D3),.enable_dir(B0_D3));   bidir_switch SK4(.port1(B1),.port2(D3),.enable_dir(B1_D3));   bidir_switch SL4(.port1(B2),.port2(D3),.enable_dir(B2_D3));   bidir_switch SM4(.port1(B3),.port2(D3),.enable_dir(B3_D3));

bidir_switch SJ5(.port1(B0),.port2(D4),.enable_dir(B0_D4));   bidir_switch SK5(.port1(B1),.port2(D4),.enable_dir(B1_D4));   bidir_switch SL5(.port1(B2),.port2(D4),.enable_dir(B2_D4));   bidir_switch SM5(.port1(B3),.port2(D4),.enable_dir(B3_D4));

bidir_switch SJ6(.port1(B0),.port2(D5),.enable_dir(B0_D5));   bidir_switch SK6(.port1(B1),.port2(D5),.enable_dir(B1_D5));   bidir_switch SL6(.port1(B2),.port2(D5),.enable_dir(B2_D5));   bidir_switch SM6(.port1(B3),.port2(D5),.enable_dir(B3_D5));

bidir_switch SJ7(.port1(B0),.port2(D6),.enable_dir(B0_D6));   bidir_switch SK7(.port1(B1),.port2(D6),.enable_dir(B1_D6));   bidir_switch SL7(.port1(B2),.port2(D6),.enable_dir(B2_D6));   bidir_switch SM7(.port1(B3),.port2(D6),.enable_dir(B3_D6));

bidir_switch SJ8(.port1(B0),.port2(D7),.enable_dir(B0_D7));   bidir_switch SK8(.port1(B1),.port2(D7),.enable_dir(B1_D7));   bidir_switch SL8(.port1(B2),.port2(D7),.enable_dir(B2_D7));   bidir_switch SM8(.port1(B3),.port2(D7),.enable_dir(B3_D7));

bidir_switch SJ9(.port1(B0),.port2(C0),.enable_dir(B0_C0));   bidir_switch SK9(.port1(B1),.port2(C0),.enable_dir(B1_C0));   bidir_switch SL9(.port1(B2),.port2(C0),.enable_dir(B2_C0));   bidir_switch SM9(.port1(B3),.port2(C0),.enable_dir(B3_C0));

bidir_switch SJ10(.port1(B0),.port2(C1),.enable_dir(B0_C1));  bidir_switch SK10(.port1(B1),.port2(C1),.enable_dir(B1_C1));  bidir_switch SL10(.port1(B2),.port2(C1),.enable_dir(B2_C1));  bidir_switch SM10(.port1(B3),.port2(C1),.enable_dir(B3_C1));

bidir_switch SJ11(.port1(B0),.port2(C2),.enable_dir(B0_C2));  bidir_switch SK11(.port1(B1),.port2(C2),.enable_dir(B1_C2));  bidir_switch SL11(.port1(B2),.port2(C2),.enable_dir(B2_C2));  bidir_switch SM11(.port1(B3),.port2(C2),.enable_dir(B3_C2));

bidir_switch SJ12(.port1(B0),.port2(C3),.enable_dir(B0_C3));  bidir_switch SK12(.port1(B1),.port2(C3),.enable_dir(B1_C3));  bidir_switch SL12(.port1(B2),.port2(C3),.enable_dir(B2_C3));  bidir_switch SM12(.port1(B3),.port2(C3),.enable_dir(B3_C3));

bidir_switch SJ13(.port1(B0),.port2(C4),.enable_dir(B0_C4));  bidir_switch SK13(.port1(B1),.port2(C4),.enable_dir(B1_C4));  bidir_switch SL13(.port1(B2),.port2(C4),.enable_dir(B2_C4));  bidir_switch SM13(.port1(B3),.port2(C4),.enable_dir(B3_C4));

bidir_switch SJ14(.port1(B0),.port2(C5),.enable_dir(B0_C5));  bidir_switch SK14(.port1(B1),.port2(C5),.enable_dir(B1_C5));  bidir_switch SL14(.port1(B2),.port2(C5),.enable_dir(B2_C5));  bidir_switch SM14(.port1(B3),.port2(C5),.enable_dir(B3_C5));

bidir_switch SJ15(.port1(B0),.port2(C6),.enable_dir(B0_C6));  bidir_switch SK15(.port1(B1),.port2(C6),.enable_dir(B1_C6));  bidir_switch SL15(.port1(B2),.port2(C6),.enable_dir(B2_C6));  bidir_switch SM15(.port1(B3),.port2(C6),.enable_dir(B3_C6));

bidir_switch SJ16(.port1(B0),.port2(C7),.enable_dir(B0_C7));  bidir_switch SK16(.port1(B1),.port2(C7),.enable_dir(B1_C7));  bidir_switch SL16(.port1(B2),.port2(C7),.enable_dir(B2_C7));  bidir_switch SM16(.port1(B3),.port2(C7),.enable_dir(B3_C7));

                                                                                                   

                                                                                                    

                                                                                                    

bidir_switch SN1(.port1(B4),.port2(D0),.enable_dir(B4_D0));	   bidir_switch SO1(.port1(B5),.port2(D0),.enable_dir(B5_D0));   bidir_switch SP1(.port1(B6),.port2(D0),.enable_dir(B6_D0));   bidir_switch SQ1(.port1(B7),.port2(D0),.enable_dir(B7_D0));

bidir_switch SN2(.port1(B4),.port2(D1),.enable_dir(B4_D1));    bidir_switch SO2(.port1(B5),.port2(D1),.enable_dir(B5_D1));   bidir_switch SP2(.port1(B6),.port2(D1),.enable_dir(B6_D1));   bidir_switch SQ2(.port1(B7),.port2(D1),.enable_dir(B7_D1));

bidir_switch SN3(.port1(B4),.port2(D2),.enable_dir(B4_D2));    bidir_switch SO3(.port1(B5),.port2(D2),.enable_dir(B5_D2));   bidir_switch SP3(.port1(B6),.port2(D2),.enable_dir(B6_D2));   bidir_switch SQ3(.port1(B7),.port2(D2),.enable_dir(B7_D2));

bidir_switch SN4(.port1(B4),.port2(D3),.enable_dir(B4_D3));    bidir_switch SO4(.port1(B5),.port2(D3),.enable_dir(B5_D3));   bidir_switch SP4(.port1(B6),.port2(D3),.enable_dir(B6_D3));   bidir_switch SQ4(.port1(B7),.port2(D3),.enable_dir(B7_D3));

bidir_switch SN5(.port1(B4),.port2(D4),.enable_dir(B4_D4));    bidir_switch SO5(.port1(B5),.port2(D4),.enable_dir(B5_D4));   bidir_switch SP5(.port1(B6),.port2(D4),.enable_dir(B6_D4));   bidir_switch SQ5(.port1(B7),.port2(D4),.enable_dir(B7_D4));

bidir_switch SN6(.port1(B4),.port2(D5),.enable_dir(B4_D5));    bidir_switch SO6(.port1(B5),.port2(D5),.enable_dir(B5_D5));   bidir_switch SP6(.port1(B6),.port2(D5),.enable_dir(B6_D5));   bidir_switch SQ6(.port1(B7),.port2(D5),.enable_dir(B7_D5));

bidir_switch SN7(.port1(B4),.port2(D6),.enable_dir(B4_D6));    bidir_switch SO7(.port1(B5),.port2(D6),.enable_dir(B5_D6));   bidir_switch SP7(.port1(B6),.port2(D6),.enable_dir(B6_D6));   bidir_switch SQ7(.port1(B7),.port2(D6),.enable_dir(B7_D6));

bidir_switch SN8(.port1(B4),.port2(D7),.enable_dir(B4_D7));    bidir_switch SO8(.port1(B5),.port2(D7),.enable_dir(B5_D7));   bidir_switch SP8(.port1(B6),.port2(D7),.enable_dir(B6_D7));   bidir_switch SQ8(.port1(B7),.port2(D7),.enable_dir(B7_D7));

bidir_switch SN9(.port1(B4),.port2(C0),.enable_dir(B4_C0));    bidir_switch SO9(.port1(B5),.port2(C0),.enable_dir(B5_C0));   bidir_switch SP9(.port1(B6),.port2(C0),.enable_dir(B6_C0));   bidir_switch SQ9(.port1(B7),.port2(C0),.enable_dir(B7_C0));

bidir_switch SN10(.port1(B4),.port2(C1),.enable_dir(B4_C1));   bidir_switch S10(.port1(B5),.port2(C1),.enable_dir(B5_C1));   bidir_switch SP10(.port1(B6),.port2(C1),.enable_dir(B6_C1));  bidir_switch SQ10(.port1(B7),.port2(C1),.enable_dir(B7_C1));

bidir_switch SN11(.port1(B4),.port2(C2),.enable_dir(B4_C2));   bidir_switch S11(.port1(B5),.port2(C2),.enable_dir(B5_C2));   bidir_switch SP11(.port1(B6),.port2(C2),.enable_dir(B6_C2));  bidir_switch SQ11(.port1(B7),.port2(C2),.enable_dir(B7_C2));

bidir_switch SN12(.port1(B4),.port2(C3),.enable_dir(B4_C3));   bidir_switch S12(.port1(B5),.port2(C3),.enable_dir(B5_C3));   bidir_switch SP12(.port1(B6),.port2(C3),.enable_dir(B6_C3));  bidir_switch SQ12(.port1(B7),.port2(C3),.enable_dir(B7_C3));

bidir_switch SN13(.port1(B4),.port2(C4),.enable_dir(B4_C4));   bidir_switch S13(.port1(B5),.port2(C4),.enable_dir(B5_C4));   bidir_switch SP13(.port1(B6),.port2(C4),.enable_dir(B6_C4));  bidir_switch SQ13(.port1(B7),.port2(C4),.enable_dir(B7_C4));

bidir_switch SN14(.port1(B4),.port2(C5),.enable_dir(B4_C5));   bidir_switch S14(.port1(B5),.port2(C5),.enable_dir(B5_C5));   bidir_switch SP14(.port1(B6),.port2(C5),.enable_dir(B6_C5));  bidir_switch SQ14(.port1(B7),.port2(C5),.enable_dir(B7_C5));

bidir_switch SN15(.port1(B4),.port2(C6),.enable_dir(B4_C6));   bidir_switch S15(.port1(B5),.port2(C6),.enable_dir(B5_C6));   bidir_switch SP15(.port1(B6),.port2(C6),.enable_dir(B6_C6));  bidir_switch SQ15(.port1(B7),.port2(C6),.enable_dir(B7_C6));

bidir_switch SN16(.port1(B4),.port2(C7),.enable_dir(B4_C7));   bidir_switch S16(.port1(B5),.port2(C7),.enable_dir(B5_C7));   bidir_switch SP16(.port1(B6),.port2(C7),.enable_dir(B6_C7));  bidir_switch SQ16(.port1(B7),.port2(C7),.enable_dir(B7_C7));

                                                                                                   

bidir_switch SR1(.port1(C0),.port2(D0),.enable_dir(C0_D0));	  bidir_switch SS1(.port1(C1),.port2(D0),.enable_dir(C1_D0));   bidir_switch ST1(.port1(C2),.port2(D0),.enable_dir(C2_D0));   bidir_switch SU1(.port1(C3),.port2(D0),.enable_dir(C3_D0));

bidir_switch SR2(.port1(C0),.port2(D1),.enable_dir(C0_D1));   bidir_switch SS2(.port1(C1),.port2(D1),.enable_dir(C1_D1));   bidir_switch ST2(.port1(C2),.port2(D1),.enable_dir(C2_D1));   bidir_switch SU2(.port1(C3),.port2(D1),.enable_dir(C3_D1));

bidir_switch SR3(.port1(C0),.port2(D2),.enable_dir(C0_D2));   bidir_switch SS3(.port1(C1),.port2(D2),.enable_dir(C1_D2));   bidir_switch ST3(.port1(C2),.port2(D2),.enable_dir(C2_D2));   bidir_switch SU3(.port1(C3),.port2(D2),.enable_dir(C3_D2));

bidir_switch SR4(.port1(C0),.port2(D3),.enable_dir(C0_D3));   bidir_switch SS4(.port1(C1),.port2(D3),.enable_dir(C1_D3));   bidir_switch ST4(.port1(C2),.port2(D3),.enable_dir(C2_D3));   bidir_switch SU4(.port1(C3),.port2(D3),.enable_dir(C3_D3));

bidir_switch SR5(.port1(C0),.port2(D4),.enable_dir(C0_D4));   bidir_switch SS5(.port1(C1),.port2(D4),.enable_dir(C1_D4));   bidir_switch ST5(.port1(C2),.port2(D4),.enable_dir(C2_D4));   bidir_switch SU5(.port1(C3),.port2(D4),.enable_dir(C3_D4));

bidir_switch SR6(.port1(C0),.port2(D5),.enable_dir(C0_D5));   bidir_switch SS6(.port1(C1),.port2(D5),.enable_dir(C1_D5));   bidir_switch ST6(.port1(C2),.port2(D5),.enable_dir(C2_D5));   bidir_switch SU6(.port1(C3),.port2(D5),.enable_dir(C3_D5));

bidir_switch SR7(.port1(C0),.port2(D6),.enable_dir(C0_D6));   bidir_switch SS7(.port1(C1),.port2(D6),.enable_dir(C1_D6));   bidir_switch ST7(.port1(C2),.port2(D6),.enable_dir(C2_D6));   bidir_switch SU7(.port1(C3),.port2(D6),.enable_dir(C3_D6));

bidir_switch SR8(.port1(C0),.port2(D7),.enable_dir(C0_D7));   bidir_switch SS8(.port1(C1),.port2(D7),.enable_dir(C1_D7));   bidir_switch ST8(.port1(C2),.port2(D7),.enable_dir(C2_D7));   bidir_switch SU8(.port1(C3),.port2(D7),.enable_dir(C3_D7));

                                                                                                    

bidir_switch SV1(.port1(C4),.port2(D0),.enable_dir(C4_D0));	  bidir_switch SW1(.port1(C5),.port2(D0),.enable_dir(C5_D0));   bidir_switch SX1(.port1(C6),.port2(D0),.enable_dir(C6_D0));   bidir_switch SY1(.port1(C7),.port2(D0),.enable_dir(C7_D0));

bidir_switch SV2(.port1(C4),.port2(D1),.enable_dir(C4_D1));   bidir_switch SW2(.port1(C5),.port2(D1),.enable_dir(C5_D1));   bidir_switch SX2(.port1(C6),.port2(D1),.enable_dir(C6_D1));   bidir_switch SY2(.port1(C7),.port2(D1),.enable_dir(C7_D1));

bidir_switch SV3(.port1(C4),.port2(D2),.enable_dir(C4_D2));   bidir_switch SW3(.port1(C5),.port2(D2),.enable_dir(C5_D2));   bidir_switch SX3(.port1(C6),.port2(D2),.enable_dir(C6_D2));   bidir_switch SY3(.port1(C7),.port2(D2),.enable_dir(C7_D2));

bidir_switch SV4(.port1(C4),.port2(D3),.enable_dir(C4_D3));   bidir_switch SW4(.port1(C5),.port2(D3),.enable_dir(C5_D3));   bidir_switch SX4(.port1(C6),.port2(D3),.enable_dir(C6_D3));   bidir_switch SY4(.port1(C7),.port2(D3),.enable_dir(C7_D3));

bidir_switch SV5(.port1(C4),.port2(D4),.enable_dir(C4_D4));   bidir_switch SW5(.port1(C5),.port2(D4),.enable_dir(C5_D4));   bidir_switch SX5(.port1(C6),.port2(D4),.enable_dir(C6_D4));   bidir_switch SY5(.port1(C7),.port2(D4),.enable_dir(C7_D4));

bidir_switch SV6(.port1(C4),.port2(D5),.enable_dir(C4_D5));   bidir_switch SW6(.port1(C5),.port2(D5),.enable_dir(C5_D5));   bidir_switch SX6(.port1(C6),.port2(D5),.enable_dir(C6_D5));   bidir_switch SY6(.port1(C7),.port2(D5),.enable_dir(C7_D5));

bidir_switch SV7(.port1(C4),.port2(D6),.enable_dir(C4_D6));   bidir_switch SW7(.port1(C5),.port2(D6),.enable_dir(C5_D6));   bidir_switch SX7(.port1(C6),.port2(D6),.enable_dir(C6_D6));   bidir_switch SY7(.port1(C7),.port2(D6),.enable_dir(C7_D6));

bidir_switch SV8(.port1(C4),.port2(D7),.enable_dir(C4_D7));   bidir_switch SW8(.port1(C5),.port2(D7),.enable_dir(C5_D7));   bidir_switch SX8(.port1(C6),.port2(D7),.enable_dir(C6_D7));   bidir_switch SY8(.port1(C7),.port2(D7),.enable_dir(C7_D7));  



`else

wire A0_B0,A0_B1,A0_B2,A0_B3,A0_B4,A0_B5,A0_B6,A0_B7,A0_C0,A0_C1,A0_C2,A0_C3,A0_C4,A0_C5,A0_C6,A0_C7,A0_D0,A0_D1,A0_D2,A0_D3,A0_D4,A0_D5,A0_D6,A0_D7,A1_B0,
A1_B1,A1_B2,A1_B3,A1_B4,A1_B5,A1_B6,A1_B7,A1_C0,A1_C1,A1_C2,A1_C3,A1_C4,A1_C5,A1_C6,A1_C7,A1_D0,A1_D1,A1_D2,A1_D3,A1_D4,A1_D5,A1_D6,A1_D7,A2_B0,A2_B1,
A2_B2,A2_B3,A2_B4,A2_B5,A2_B6,A2_B7,A2_C0,A2_C1,A2_C2,A2_C3,A2_C4,A2_C5,A2_C6,A2_C7,A2_D0,A2_D1,A2_D2,A2_D3,A2_D4,A2_D5,A2_D6,A2_D7,A3_B0,A3_B1,A3_B2,
A3_B3,A3_B4,A3_B5,A3_B6,A3_B7,A3_C0,A3_C1,A3_C2,A3_C3,A3_C4,A3_C5,A3_C6,A3_C7,A3_D0,A3_D1,A3_D2,A3_D3,A3_D4,A3_D5,A3_D6,A3_D7,A4_B0,A4_B1,A4_B2,A4_B3,
A4_B4,A4_B5,A4_B6,A4_B7,A4_C0,A4_C1,A4_C2,A4_C3,A4_C4,A4_C5,A4_C6,A4_C7,A4_D0,A4_D1,A4_D2,A4_D3,A4_D4,A4_D5,A4_D6,A4_D7,A5_B0,A5_B1,A5_B2,A5_B3,A5_B4,
A5_B5,A5_B6,A5_B7,A5_C0,A5_C1,A5_C2,A5_C3,A5_C4,A5_C5,A5_C6,A5_C7,A5_D0,A5_D1,A5_D2,A5_D3,A5_D4,A5_D5,A5_D6,A5_D7,A6_B0,A6_B1,A6_B2,A6_B3,A6_B4,A6_B5,
A6_B6,A6_B7,A6_C0,A6_C1,A6_C2,A6_C3,A6_C4,A6_C5,A6_C6,A6_C7,A6_D0,A6_D1,A6_D2,A6_D3,A6_D4,A6_D5,A6_D6,A6_D7,A7_B0,A7_B1,A7_B2,A7_B3,A7_B4,A7_B5,A7_B6,
A7_B7,A7_C0,A7_C1,A7_C2,A7_C3,A7_C4,A7_C5,A7_C6,A7_C7,A7_D0,A7_D1,A7_D2,A7_D3,A7_D4,A7_D5,A7_D6,A7_D7,B0_D0,B0_D1,B0_D2,B0_D3,B0_D4,B0_D5,B0_D6,B0_D7,
B0_C0,B0_C1,B0_C2,B0_C3,B0_C4,B0_C5,B0_C6,B0_C7,B1_D0,B1_D1,B1_D2,B1_D3,B1_D4,B1_D5,B1_D6,B1_D7,B1_C0,B1_C1,B1_C2,B1_C3,B1_C4,B1_C5,B1_C6,B1_C7,B2_D0,
B2_D1,B2_D2,B2_D3,B2_D4,B2_D5,B2_D6,B2_D7,B2_C0,B2_C1,B2_C2,B2_C3,B2_C4,B2_C5,B2_C6,B2_C7,B3_D0,B3_D1,B3_D2,B3_D3,B3_D4,B3_D5,B3_D6,B3_D7,B3_C0,B3_C1,
B3_C2,B3_C3,B3_C4,B3_C5,B3_C6,B3_C7,B4_D0,B4_D1,B4_D2,B4_D3,B4_D4,B4_D5,B4_D6,B4_D7,B4_C0,B4_C1,B4_C2,B4_C3,B4_C4,B4_C5,B4_C6,B4_C7,B5_D0,B5_D1,B5_D2,
B5_D3,B5_D4,B5_D5,B5_D6,B5_D7,B5_C0,B5_C1,B5_C2,B5_C3,B5_C4,B5_C5,B5_C6,B5_C7,B6_D0,B6_D1,B6_D2,B6_D3,B6_D4,B6_D5,B6_D6,B6_D7,B6_C0,B6_C1,B6_C2,B6_C3,
B6_C4,B6_C5,B6_C6,B6_C7,B7_D0,B7_D1,B7_D2,B7_D3,B7_D4,B7_D5,B7_D6,B7_D7,B7_C0,B7_C1,B7_C2,B7_C3,B7_C4,B7_C5,B7_C6,B7_C7,C0_D0,C0_D1,C0_D2,C0_D3,C0_D4,
C0_D5,C0_D6,C0_D7,C1_D0,C1_D1,C1_D2,C1_D3,C1_D4,C1_D5,C1_D6,C1_D7,C2_D0,C2_D1,C2_D2,C2_D3,C2_D4,C2_D5,C2_D6,C2_D7,C3_D0,C3_D1,C3_D2,C3_D3,C3_D4,C3_D5,
C3_D6,C3_D7,C4_D0,C4_D1,C4_D2,C4_D3,C4_D4,C4_D5,C4_D6,C4_D7,C5_D0,C5_D1,C5_D2,C5_D3,C5_D4,C5_D5,C5_D6,C5_D7,C6_D0,C6_D1,C6_D2,C6_D3,C6_D4,C6_D5,C6_D6,
C6_D7,C7_D0,C7_D1,C7_D2,C7_D3,C7_D4,C7_D5,C7_D6,C7_D7;

switch_block_config Bidir_switch (.bit_in(bit_in),.bit_out(bit_out),.prgm_b(prgm_b),.sb_prgm_b(sb_prgm_b),.clk(clk),.reset(reset),
.A0_B0(A0_B0),.A0_B1(A0_B1),.A0_B2(A0_B2),.A0_B3(A0_B3),.A0_B4(A0_B4),.A0_B5(A0_B5),.A0_B6(A0_B6),.A0_B7(A0_B7),.A0_C0(A0_C0),.A0_C1(A0_C1),.A0_C2(A0_C2),.A0_C3(A0_C3),.A0_C4(A0_C4),.A0_C5(A0_C5),.A0_C6(A0_C6),.A0_C7(A0_C7),.A0_D0(A0_D0),.A0_D1(A0_D1),.A0_D2(A0_D2),.A0_D3(A0_D3),.A0_D4(A0_D4),.A0_D5(A0_D5),.A0_D6(A0_D6),.A0_D7(A0_D7),.A1_B0(A1_B0),
.A1_B1(A1_B1),.A1_B2(A1_B2),.A1_B3(A1_B3),.A1_B4(A1_B4),.A1_B5(A1_B5),.A1_B6(A1_B6),.A1_B7(A1_B7),.A1_C0(A1_C0),.A1_C1(A1_C1),.A1_C2(A1_C2),.A1_C3(A1_C3),.A1_C4(A1_C4),.A1_C5(A1_C5),.A1_C6(A1_C6),.A1_C7(A1_C7),.A1_D0(A1_D0),.A1_D1(A1_D1),.A1_D2(A1_D2),.A1_D3(A1_D3),.A1_D4(A1_D4),.A1_D5(A1_D5),.A1_D6(A1_D6),.A1_D7(A1_D7),.A2_B0(A2_B0),.A2_B1(A2_B1),
.A2_B2(A2_B2),.A2_B3(A2_B3),.A2_B4(A2_B4),.A2_B5(A2_B5),.A2_B6(A2_B6),.A2_B7(A2_B7),.A2_C0(A2_C0),.A2_C1(A2_C1),.A2_C2(A2_C2),.A2_C3(A2_C3),.A2_C4(A2_C4),.A2_C5(A2_C5),.A2_C6(A2_C6),.A2_C7(A2_C7),.A2_D0(A2_D0),.A2_D1(A2_D1),.A2_D2(A2_D2),.A2_D3(A2_D3),.A2_D4(A2_D4),.A2_D5(A2_D5),.A2_D6(A2_D6),.A2_D7(A2_D7),.A3_B0(A3_B0),.A3_B1(A3_B1),.A3_B2(A3_B2),
.A3_B3(A3_B3),.A3_B4(A3_B4),.A3_B5(A3_B5),.A3_B6(A3_B6),.A3_B7(A3_B7),.A3_C0(A3_C0),.A3_C1(A3_C1),.A3_C2(A3_C2),.A3_C3(A3_C3),.A3_C4(A3_C4),.A3_C5(A3_C5),.A3_C6(A3_C6),.A3_C7(A3_C7),.A3_D0(A3_D0),.A3_D1(A3_D1),.A3_D2(A3_D2),.A3_D3(A3_D3),.A3_D4(A3_D4),.A3_D5(A3_D5),.A3_D6(A3_D6),.A3_D7(A3_D7),.A4_B0(A4_B0),.A4_B1(A4_B1),.A4_B2(A4_B2),.A4_B3(A4_B3),
.A4_B4(A4_B4),.A4_B5(A4_B5),.A4_B6(A4_B6),.A4_B7(A4_B7),.A4_C0(A4_C0),.A4_C1(A4_C1),.A4_C2(A4_C2),.A4_C3(A4_C3),.A4_C4(A4_C4),.A4_C5(A4_C5),.A4_C6(A4_C6),.A4_C7(A4_C7),.A4_D0(A4_D0),.A4_D1(A4_D1),.A4_D2(A4_D2),.A4_D3(A4_D3),.A4_D4(A4_D4),.A4_D5(A4_D5),.A4_D6(A4_D6),.A4_D7(A4_D7),.A5_B0(A5_B0),.A5_B1(A5_B1),.A5_B2(A5_B2),.A5_B3(A5_B3),.A5_B4(A5_B4),
.A5_B5(A5_B5),.A5_B6(A5_B6),.A5_B7(A5_B7),.A5_C0(A5_C0),.A5_C1(A5_C1),.A5_C2(A5_C2),.A5_C3(A5_C3),.A5_C4(A5_C4),.A5_C5(A5_C5),.A5_C6(A5_C6),.A5_C7(A5_C7),.A5_D0(A5_D0),.A5_D1(A5_D1),.A5_D2(A5_D2),.A5_D3(A5_D3),.A5_D4(A5_D4),.A5_D5(A5_D5),.A5_D6(A5_D6),.A5_D7(A5_D7),.A6_B0(A6_B0),.A6_B1(A6_B1),.A6_B2(A6_B2),.A6_B3(A6_B3),.A6_B4(A6_B4),.A6_B5(A6_B5),
.A6_B6(A6_B6),.A6_B7(A6_B7),.A6_C0(A6_C0),.A6_C1(A6_C1),.A6_C2(A6_C2),.A6_C3(A6_C3),.A6_C4(A6_C4),.A6_C5(A6_C5),.A6_C6(A6_C6),.A6_C7(A6_C7),.A6_D0(A6_D0),.A6_D1(A6_D1),.A6_D2(A6_D2),.A6_D3(A6_D3),.A6_D4(A6_D4),.A6_D5(A6_D5),.A6_D6(A6_D6),.A6_D7(A6_D7),.A7_B0(A7_B0),.A7_B1(A7_B1),.A7_B2(A7_B2),.A7_B3(A7_B3),.A7_B4(A7_B4),.A7_B5(A7_B5),.A7_B6(A7_B6),
.A7_B7(A7_B7),.A7_C0(A7_C0),.A7_C1(A7_C1),.A7_C2(A7_C2),.A7_C3(A7_C3),.A7_C4(A7_C4),.A7_C5(A7_C5),.A7_C6(A7_C6),.A7_C7(A7_C7),.A7_D0(A7_D0),.A7_D1(A7_D1),.A7_D2(A7_D2),.A7_D3(A7_D3),.A7_D4(A7_D4),.A7_D5(A7_D5),.A7_D6(A7_D6),.A7_D7(A7_D7),.B0_D0(B0_D0),.B0_D1(B0_D1),.B0_D2(B0_D2),.B0_D3(B0_D3),.B0_D4(B0_D4),.B0_D5(B0_D5),.B0_D6(B0_D6),.B0_D7(B0_D7),
.B0_C0(B0_C0),.B0_C1(B0_C1),.B0_C2(B0_C2),.B0_C3(B0_C3),.B0_C4(B0_C4),.B0_C5(B0_C5),.B0_C6(B0_C6),.B0_C7(B0_C7),.B1_D0(B1_D0),.B1_D1(B1_D1),.B1_D2(B1_D2),.B1_D3(B1_D3),.B1_D4(B1_D4),.B1_D5(B1_D5),.B1_D6(B1_D6),.B1_D7(B1_D7),.B1_C0(B1_C0),.B1_C1(B1_C1),.B1_C2(B1_C2),.B1_C3(B1_C3),.B1_C4(B1_C4),.B1_C5(B1_C5),.B1_C6(B1_C6),.B1_C7(B1_C7),.B2_D0(B2_D0),
.B2_D1(B2_D1),.B2_D2(B2_D2),.B2_D3(B2_D3),.B2_D4(B2_D4),.B2_D5(B2_D5),.B2_D6(B2_D6),.B2_D7(B2_D7),.B2_C0(B2_C0),.B2_C1(B2_C1),.B2_C2(B2_C2),.B2_C3(B2_C3),.B2_C4(B2_C4),.B2_C5(B2_C5),.B2_C6(B2_C6),.B2_C7(B2_C7),.B3_D0(B3_D0),.B3_D1(B3_D1),.B3_D2(B3_D2),.B3_D3(B3_D3),.B3_D4(B3_D4),.B3_D5(B3_D5),.B3_D6(B3_D6),.B3_D7(B3_D7),.B3_C0(B3_C0),.B3_C1(B3_C1),
.B3_C2(B3_C2),.B3_C3(B3_C3),.B3_C4(B3_C4),.B3_C5(B3_C5),.B3_C6(B3_C6),.B3_C7(B3_C7),.B4_D0(B4_D0),.B4_D1(B4_D1),.B4_D2(B4_D2),.B4_D3(B4_D3),.B4_D4(B4_D4),.B4_D5(B4_D5),.B4_D6(B4_D6),.B4_D7(B4_D7),.B4_C0(B4_C0),.B4_C1(B4_C1),.B4_C2(B4_C2),.B4_C3(B4_C3),.B4_C4(B4_C4),.B4_C5(B4_C5),.B4_C6(B4_C6),.B4_C7(B4_C7),.B5_D0(B5_D0),.B5_D1(B5_D1),.B5_D2(B5_D2),
.B5_D3(B5_D3),.B5_D4(B5_D4),.B5_D5(B5_D5),.B5_D6(B5_D6),.B5_D7(B5_D7),.B5_C0(B5_C0),.B5_C1(B5_C1),.B5_C2(B5_C2),.B5_C3(B5_C3),.B5_C4(B5_C4),.B5_C5(B5_C5),.B5_C6(B5_C6),.B5_C7(B5_C7),.B6_D0(B6_D0),.B6_D1(B6_D1),.B6_D2(B6_D2),.B6_D3(B6_D3),.B6_D4(B6_D4),.B6_D5(B6_D5),.B6_D6(B6_D6),.B6_D7(B6_D7),.B6_C0(B6_C0),.B6_C1(B6_C1),.B6_C2(B6_C2),.B6_C3(B6_C3),
.B6_C4(B6_C4),.B6_C5(B6_C5),.B6_C6(B6_C6),.B6_C7(B6_C7),.B7_D0(B7_D0),.B7_D1(B7_D1),.B7_D2(B7_D2),.B7_D3(B7_D3),.B7_D4(B7_D4),.B7_D5(B7_D5),.B7_D6(B7_D6),.B7_D7(B7_D7),.B7_C0(B7_C0),.B7_C1(B7_C1),.B7_C2(B7_C2),.B7_C3(B7_C3),.B7_C4(B7_C4),.B7_C5(B7_C5),.B7_C6(B7_C6),.B7_C7(B7_C7),.C0_D0(C0_D0),.C0_D1(C0_D1),.C0_D2(C0_D2),.C0_D3(C0_D3),.C0_D4(C0_D4),
.C0_D5(C0_D5),.C0_D6(C0_D6),.C0_D7(C0_D7),.C1_D0(C1_D0),.C1_D1(C1_D1),.C1_D2(C1_D2),.C1_D3(C1_D3),.C1_D4(C1_D4),.C1_D5(C1_D5),.C1_D6(C1_D6),.C1_D7(C1_D7),.C2_D0(C2_D0),.C2_D1(C2_D1),.C2_D2(C2_D2),.C2_D3(C2_D3),.C2_D4(C2_D4),.C2_D5(C2_D5),.C2_D6(C2_D6),.C2_D7(C2_D7),.C3_D0(C3_D0),.C3_D1(C3_D1),.C3_D2(C3_D2),.C3_D3(C3_D3),.C3_D4(C3_D4),.C3_D5(C3_D5),
.C3_D6(C3_D6),.C3_D7(C3_D7),.C4_D0(C4_D0),.C4_D1(C4_D1),.C4_D2(C4_D2),.C4_D3(C4_D3),.C4_D4(C4_D4),.C4_D5(C4_D5),.C4_D6(C4_D6),.C4_D7(C4_D7),.C5_D0(C5_D0),.C5_D1(C5_D1),.C5_D2(C5_D2),.C5_D3(C5_D3),.C5_D4(C5_D4),.C5_D5(C5_D5),.C5_D6(C5_D6),.C5_D7(C5_D7),.C6_D0(C6_D0),.C6_D1(C6_D1),.C6_D2(C6_D2),.C6_D3(C6_D3),.C6_D4(C6_D4),.C6_D5(C6_D5),.C6_D6(C6_D6),
.C6_D7(C6_D7),.C7_D0(C7_D0),.C7_D1(C7_D1),.C7_D2(C7_D2),.C7_D3(C7_D3),.C7_D4(C7_D4),.C7_D5(C7_D5),.C7_D6(C7_D6),.C7_D7(C7_D7));

tranif1(B0,A0,A0_B0);	tranif1(B0,A1,A1_B0);   tranif1(B0,A2,A2_B0);	tranif1(B0,A3,A3_B0);
tranif1(B1,A0,A0_B1);   tranif1(B1,A1,A1_B1);   tranif1(B1,A2,A2_B1);   tranif1(B1,A3,A3_B1);
tranif1(B2,A0,A0_B2);   tranif1(B2,A1,A1_B2);   tranif1(B2,A2,A2_B2);   tranif1(B2,A3,A3_B2);
tranif1(B3,A0,A0_B3);   tranif1(B3,A1,A1_B3);   tranif1(B3,A2,A2_B3);   tranif1(B3,A3,A3_B3);
tranif1(B4,A0,A0_B4);   tranif1(B4,A1,A1_B4);   tranif1(B4,A2,A2_B4);   tranif1(B4,A3,A3_B4);
tranif1(B5,A0,A0_B5);   tranif1(B5,A1,A1_B5);   tranif1(B5,A2,A2_B5);   tranif1(B5,A3,A3_B5);
tranif1(B6,A0,A0_B6);   tranif1(B6,A1,A1_B6);   tranif1(B6,A2,A2_B6);   tranif1(B6,A3,A3_B6);
tranif1(B7,A0,A0_B7);   tranif1(B7,A1,A1_B7);   tranif1(B7,A2,A2_B7);   tranif1(B7,A3,A3_B7);
tranif1(C0,A0,A0_C0);   tranif1(C0,A1,A1_C0);   tranif1(C0,A2,A2_C0);   tranif1(C0,A3,A3_C0);
tranif1(C1,A0,A0_C1);   tranif1(C1,A1,A1_C1);   tranif1(C1,A2,A2_C1);   tranif1(C1,A3,A3_C1);
tranif1(C2,A0,A0_C2);   tranif1(C2,A1,A1_C2);   tranif1(C2,A2,A2_C2);   tranif1(C2,A3,A3_C2);
tranif1(C3,A0,A0_C3);   tranif1(C3,A1,A1_C3);   tranif1(C3,A2,A2_C3);   tranif1(C3,A3,A3_C3);
tranif1(C4,A0,A0_C4);   tranif1(C4,A1,A1_C4);   tranif1(C4,A2,A2_C4);   tranif1(C4,A3,A3_C4);
tranif1(C5,A0,A0_C5);   tranif1(C5,A1,A1_C5);   tranif1(C5,A2,A2_C5);   tranif1(C5,A3,A3_C5);
tranif1(C6,A0,A0_C6);   tranif1(C6,A1,A1_C6);   tranif1(C6,A2,A2_C6);   tranif1(C6,A3,A3_C6);
tranif1(C7,A0,A0_C7);   tranif1(C7,A1,A1_C7);   tranif1(C7,A2,A2_C7);   tranif1(C7,A3,A3_C7);
tranif1(D0,A0,A0_D0);   tranif1(D0,A1,A1_D0);   tranif1(D0,A2,A2_D0);   tranif1(D0,A3,A3_D0);
tranif1(D1,A0,A0_D1);   tranif1(D1,A1,A1_D1);   tranif1(D1,A2,A2_D1);   tranif1(D1,A3,A3_D1);
tranif1(D2,A0,A0_D2);   tranif1(D2,A1,A1_D2);   tranif1(D2,A2,A2_D2);   tranif1(D2,A3,A3_D2);
tranif1(D3,A0,A0_D3);   tranif1(D3,A1,A1_D3);   tranif1(D3,A2,A2_D3);   tranif1(D3,A3,A3_D3);
tranif1(D4,A0,A0_D4);   tranif1(D4,A1,A1_D4);   tranif1(D4,A2,A2_D4);   tranif1(D4,A3,A3_D4);
tranif1(D5,A0,A0_D5);   tranif1(D5,A1,A1_D5);   tranif1(D5,A2,A2_D5);   tranif1(D5,A3,A3_D5);
tranif1(D6,A0,A0_D6);   tranif1(D6,A1,A1_D6);   tranif1(D6,A2,A2_D6);   tranif1(D6,A3,A3_D6);
tranif1(D7,A0,A0_D7);   tranif1(D7,A1,A1_D7);   tranif1(D7,A2,A2_D7);   tranif1(D7,A3,A3_D7);



tranif1(B0,A4,A4_B0);	tranif1(B0,A5,A5_B0);   tranif1(B0,A6,A6_B0);	tranif1(B0,A7,A7_B0);
tranif1(B1,A4,A4_B1);   tranif1(B1,A5,A5_B1);   tranif1(B1,A6,A6_B1);   tranif1(B1,A7,A7_B1);
tranif1(B2,A4,A4_B2);   tranif1(B2,A5,A5_B2);   tranif1(B2,A6,A6_B2);   tranif1(B2,A7,A7_B2);
tranif1(B3,A4,A4_B3);   tranif1(B3,A5,A5_B3);   tranif1(B3,A6,A6_B3);   tranif1(B3,A7,A7_B3);
tranif1(B4,A4,A4_B4);   tranif1(B4,A5,A5_B4);   tranif1(B4,A6,A6_B4);   tranif1(B4,A7,A7_B4);
tranif1(B5,A4,A4_B5);   tranif1(B5,A5,A5_B5);   tranif1(B5,A6,A6_B5);   tranif1(B5,A7,A7_B5);
tranif1(B6,A4,A4_B6);   tranif1(B6,A5,A5_B6);   tranif1(B6,A6,A6_B6);   tranif1(B6,A7,A7_B6);
tranif1(B7,A4,A4_B7);   tranif1(B7,A5,A5_B7);   tranif1(B7,A6,A6_B7);   tranif1(B7,A7,A7_B7);
tranif1(C0,A4,A4_C0);   tranif1(C0,A5,A5_C0);   tranif1(C0,A6,A6_C0);   tranif1(C0,A7,A7_C0);
tranif1(C1,A4,A4_C1);   tranif1(C1,A5,A5_C1);   tranif1(C1,A6,A6_C1);   tranif1(C1,A7,A7_C1);
tranif1(C2,A4,A4_C2);   tranif1(C2,A5,A5_C2);   tranif1(C2,A6,A6_C2);   tranif1(C2,A7,A7_C2);
tranif1(C3,A4,A4_C3);   tranif1(C3,A5,A5_C3);   tranif1(C3,A6,A6_C3);   tranif1(C3,A7,A7_C3);
tranif1(C4,A4,A4_C4);   tranif1(C4,A5,A5_C4);   tranif1(C4,A6,A6_C4);   tranif1(C4,A7,A7_C4);
tranif1(C5,A4,A4_C5);   tranif1(C5,A5,A5_C5);   tranif1(C5,A6,A6_C5);   tranif1(C5,A7,A7_C5);
tranif1(C6,A4,A4_C6);   tranif1(C6,A5,A5_C6);   tranif1(C6,A6,A6_C6);   tranif1(C6,A7,A7_C6);
tranif1(C7,A4,A4_C7);   tranif1(C7,A5,A5_C7);   tranif1(C7,A6,A6_C7);   tranif1(C7,A7,A7_C7);
tranif1(D0,A4,A4_D0);   tranif1(D0,A5,A5_D0);   tranif1(D0,A6,A6_D0);   tranif1(D0,A7,A7_D0);
tranif1(D1,A4,A4_D1);   tranif1(D1,A5,A5_D1);   tranif1(D1,A6,A6_D1);   tranif1(D1,A7,A7_D1);
tranif1(D2,A4,A4_D2);   tranif1(D2,A5,A5_D2);   tranif1(D2,A6,A6_D2);   tranif1(D2,A7,A7_D2);
tranif1(D3,A4,A4_D3);   tranif1(D3,A5,A5_D3);   tranif1(D3,A6,A6_D3);   tranif1(D3,A7,A7_D3);
tranif1(D4,A4,A4_D4);   tranif1(D4,A5,A5_D4);   tranif1(D4,A6,A6_D4);   tranif1(D4,A7,A7_D4);
tranif1(D5,A4,A4_D5);   tranif1(D5,A5,A5_D5);   tranif1(D5,A6,A6_D5);   tranif1(D5,A7,A7_D5);
tranif1(D6,A4,A4_D6);   tranif1(D6,A5,A5_D6);   tranif1(D6,A6,A6_D6);   tranif1(D6,A7,A7_D6);
tranif1(D7,A4,A4_D7);   tranif1(D7,A5,A5_D7);   tranif1(D7,A6,A6_D7);   tranif1(D7,A7,A7_D7);


tranif1(D0,B0,B0_D0);	tranif1(D0,B1,B1_D0);   tranif1(D0,B2,B2_D0);	tranif1(D0,B3,B3_D0);
tranif1(D1,B0,B0_D1);   tranif1(D1,B1,B1_D1);   tranif1(D1,B2,B2_D1);   tranif1(D1,B3,B3_D1);
tranif1(D2,B0,B0_D2);   tranif1(D2,B1,B1_D2);   tranif1(D2,B2,B2_D2);   tranif1(D2,B3,B3_D2);
tranif1(D3,B0,B0_D3);   tranif1(D3,B1,B1_D3);   tranif1(D3,B2,B2_D3);   tranif1(D3,B3,B3_D3);
tranif1(D4,B0,B0_D4);   tranif1(D4,B1,B1_D4);   tranif1(D4,B2,B2_D4);   tranif1(D4,B3,B3_D4);
tranif1(D5,B0,B0_D5);   tranif1(D5,B1,B1_D5);   tranif1(D5,B2,B2_D5);   tranif1(D5,B3,B3_D5);
tranif1(D6,B0,B0_D6);   tranif1(D6,B1,B1_D6);   tranif1(D6,B2,B2_D6);   tranif1(D6,B3,B3_D6);
tranif1(D7,B0,B0_D7);   tranif1(D7,B1,B1_D7);   tranif1(D7,B2,B2_D7);   tranif1(D7,B3,B3_D7);
tranif1(C0,B0,B0_C0);   tranif1(C0,B1,B1_C0);   tranif1(C0,B2,B2_C0);   tranif1(C0,B3,B3_C0);
tranif1(C1,B0,B0_C1);   tranif1(C1,B1,B1_C1);   tranif1(C1,B2,B2_C1);   tranif1(C1,B3,B3_C1);
tranif1(C2,B0,B0_C2);   tranif1(C2,B1,B1_C2);   tranif1(C2,B2,B2_C2);   tranif1(C2,B3,B3_C2);
tranif1(C3,B0,B0_C3);   tranif1(C3,B1,B1_C3);   tranif1(C3,B2,B2_C3);   tranif1(C3,B3,B3_C3);
tranif1(C4,B0,B0_C4);   tranif1(C4,B1,B1_C4);   tranif1(C4,B2,B2_C4);   tranif1(C4,B3,B3_C4);
tranif1(C5,B0,B0_C5);   tranif1(C5,B1,B1_C5);   tranif1(C5,B2,B2_C5);   tranif1(C5,B3,B3_C5);
tranif1(C6,B0,B0_C6);   tranif1(C6,B1,B1_C6);   tranif1(C6,B2,B2_C6);   tranif1(C6,B3,B3_C6);
tranif1(C7,B0,B0_C7);   tranif1(C7,B1,B1_C7);   tranif1(C7,B2,B2_C7);   tranif1(C7,B3,B3_C7);



tranif1(D0,B4,B4_D0);	tranif1(D0,B5,B5_D0);   tranif1(D0,B6,B6_D0);	tranif1(D0,B7,B7_D0);
tranif1(D1,B4,B4_D1);   tranif1(D1,B5,B5_D1);   tranif1(D1,B6,B6_D1);   tranif1(D1,B7,B7_D1);
tranif1(D2,B4,B4_D2);   tranif1(D2,B5,B5_D2);   tranif1(D2,B6,B6_D2);   tranif1(D2,B7,B7_D2);
tranif1(D3,B4,B4_D3);   tranif1(D3,B5,B5_D3);   tranif1(D3,B6,B6_D3);   tranif1(D3,B7,B7_D3);
tranif1(D4,B4,B4_D4);   tranif1(D4,B5,B5_D4);   tranif1(D4,B6,B6_D4);   tranif1(D4,B7,B7_D4);
tranif1(D5,B4,B4_D5);   tranif1(D5,B5,B5_D5);   tranif1(D5,B6,B6_D5);   tranif1(D5,B7,B7_D5);
tranif1(D6,B4,B4_D6);   tranif1(D6,B5,B5_D6);   tranif1(D6,B6,B6_D6);   tranif1(D6,B7,B7_D6);
tranif1(D7,B4,B4_D7);   tranif1(D7,B5,B5_D7);   tranif1(D7,B6,B6_D7);   tranif1(D7,B7,B7_D7);
tranif1(C0,B4,B4_C0);   tranif1(C0,B5,B5_C0);   tranif1(C0,B6,B6_C0);   tranif1(C0,B7,B7_C0);
tranif1(C1,B4,B4_C1);   tranif1(C1,B5,B5_C1);   tranif1(C1,B6,B6_C1);   tranif1(C1,B7,B7_C1);
tranif1(C2,B4,B4_C2);   tranif1(C2,B5,B5_C2);   tranif1(C2,B6,B6_C2);   tranif1(C2,B7,B7_C2);
tranif1(C3,B4,B4_C3);   tranif1(C3,B5,B5_C3);   tranif1(C3,B6,B6_C3);   tranif1(C3,B7,B7_C3);
tranif1(C4,B4,B4_C4);   tranif1(C4,B5,B5_C4);   tranif1(C4,B6,B6_C4);   tranif1(C4,B7,B7_C4);
tranif1(C5,B4,B4_C5);   tranif1(C5,B5,B5_C5);   tranif1(C5,B6,B6_C5);   tranif1(C5,B7,B7_C5);
tranif1(C6,B4,B4_C6);   tranif1(C6,B5,B5_C6);   tranif1(C6,B6,B6_C6);   tranif1(C6,B7,B7_C6);
tranif1(C7,B4,B4_C7);   tranif1(C7,B5,B5_C7);   tranif1(C7,B6,B6_C7);   tranif1(C7,B7,B7_C7);

tranif1(D0,C0,C0_D0);	tranif1(D0,C1,C1_D0);   tranif1(D0,C2,C2_D0);	tranif1(D0,C3,C3_D0);
tranif1(D1,C0,C0_D1);   tranif1(D1,C1,C1_D1);   tranif1(D1,C2,C2_D1);   tranif1(D1,C3,C3_D1);
tranif1(D2,C0,C0_D2);   tranif1(D2,C1,C1_D2);   tranif1(D2,C2,C2_D2);   tranif1(D2,C3,C3_D2);
tranif1(D3,C0,C0_D3);   tranif1(D3,C1,C1_D3);   tranif1(D3,C2,C2_D3);   tranif1(D3,C3,C3_D3);
tranif1(D4,C0,C0_D4);   tranif1(D4,C1,C1_D4);   tranif1(D4,C2,C2_D4);   tranif1(D4,C3,C3_D4);
tranif1(D5,C0,C0_D5);   tranif1(D5,C1,C1_D5);   tranif1(D5,C2,C2_D5);   tranif1(D5,C3,C3_D5);
tranif1(D6,C0,C0_D6);   tranif1(D6,C1,C1_D6);   tranif1(D6,C2,C2_D6);   tranif1(D6,C3,C3_D6);
tranif1(D7,C0,C0_D7);   tranif1(D7,C1,C1_D7);   tranif1(D7,C2,C2_D7);   tranif1(D7,C3,C3_D7);

tranif1(D0,C4,C4_D0);	tranif1(D0,C5,C5_D0);   tranif1(D0,C6,C6_D0);	tranif1(D0,C7,C7_D0);
tranif1(D1,C4,C4_D1);   tranif1(D1,C5,C5_D1);   tranif1(D1,C6,C6_D1);   tranif1(D1,C7,C7_D1);
tranif1(D2,C4,C4_D2);   tranif1(D2,C5,C5_D2);   tranif1(D2,C6,C6_D2);   tranif1(D2,C7,C7_D2);
tranif1(D3,C4,C4_D3);   tranif1(D3,C5,C5_D3);   tranif1(D3,C6,C6_D3);   tranif1(D3,C7,C7_D3);
tranif1(D4,C4,C4_D4);   tranif1(D4,C5,C5_D4);   tranif1(D4,C6,C6_D4);   tranif1(D4,C7,C7_D4);
tranif1(D5,C4,C4_D5);   tranif1(D5,C5,C5_D5);   tranif1(D5,C6,C6_D5);   tranif1(D5,C7,C7_D5);
tranif1(D6,C4,C4_D6);   tranif1(D6,C5,C5_D6);   tranif1(D6,C6,C6_D6);   tranif1(D6,C7,C7_D6);
tranif1(D7,C4,C4_D7);   tranif1(D7,C5,C5_D7);   tranif1(D7,C6,C6_D7);   tranif1(D7,C7,C7_D7);

`endif

endmodule
